module MacUnit(
  input  [7:0]  io_in_a, // @[src/main/scala/gemmini/PE.scala 16:14]
  input  [7:0]  io_in_b, // @[src/main/scala/gemmini/PE.scala 16:14]
  input  [19:0] io_in_c, // @[src/main/scala/gemmini/PE.scala 16:14]
  output [19:0] io_out_d // @[src/main/scala/gemmini/PE.scala 16:14]
);
  wire [15:0] _io_out_d_T = $signed(io_in_a) * $signed(io_in_b); // @[src/main/scala/gemmini/Arithmetic.scala 37:49]
  wire [19:0] _GEN_0 = {{4{_io_out_d_T[15]}},_io_out_d_T}; // @[src/main/scala/gemmini/Arithmetic.scala 37:54]
  assign io_out_d = $signed(_GEN_0) + $signed(io_in_c); // @[src/main/scala/gemmini/Arithmetic.scala 37:54]
endmodule
module PE(
  input         clock,
  input  [7:0]  io_in_a, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [19:0] io_in_b, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [19:0] io_in_d, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [7:0]  io_out_a, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [19:0] io_out_b, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [19:0] io_out_c, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_control_dataflow, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_control_propagate, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [4:0]  io_in_control_shift, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_control_dataflow, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_control_propagate, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [4:0]  io_out_control_shift, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [1:0]  io_in_id, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [1:0]  io_out_id, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_last, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_last, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_valid, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_valid // @[src/main/scala/gemmini/PE.scala 35:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] mac_unit_io_in_a; // @[src/main/scala/gemmini/PE.scala 64:24]
  wire [7:0] mac_unit_io_in_b; // @[src/main/scala/gemmini/PE.scala 64:24]
  wire [19:0] mac_unit_io_in_c; // @[src/main/scala/gemmini/PE.scala 64:24]
  wire [19:0] mac_unit_io_out_d; // @[src/main/scala/gemmini/PE.scala 64:24]
  reg [7:0] c1; // @[src/main/scala/gemmini/PE.scala 70:15]
  reg [7:0] c2; // @[src/main/scala/gemmini/PE.scala 71:15]
  wire [7:0] _GEN_7 = io_in_control_propagate ? $signed(c1) : $signed(c2); // @[src/main/scala/gemmini/PE.scala 119:30 120:16 126:16]
  wire [19:0] _GEN_11 = io_in_control_propagate ? $signed(io_in_d) : $signed({{12{c1[7]}},c1}); // @[src/main/scala/gemmini/PE.scala 119:30 124:10 70:15]
  wire [19:0] _GEN_12 = io_in_control_propagate ? $signed({{12{c2[7]}},c2}) : $signed(io_in_d); // @[src/main/scala/gemmini/PE.scala 119:30 130:10 71:15]
  wire [19:0] _GEN_27 = ~io_in_valid ? $signed({{12{c1[7]}},c1}) : $signed(_GEN_11); // @[src/main/scala/gemmini/PE.scala 141:17 142:8]
  wire [19:0] _GEN_28 = ~io_in_valid ? $signed({{12{c2[7]}},c2}) : $signed(_GEN_12); // @[src/main/scala/gemmini/PE.scala 141:17 143:8]
  MacUnit mac_unit ( // @[src/main/scala/gemmini/PE.scala 64:24]
    .io_in_a(mac_unit_io_in_a),
    .io_in_b(mac_unit_io_in_b),
    .io_in_c(mac_unit_io_in_c),
    .io_out_d(mac_unit_io_out_d)
  );
  assign io_out_a = io_in_a; // @[src/main/scala/gemmini/PE.scala 79:12]
  assign io_out_b = mac_unit_io_out_d; // @[src/main/scala/gemmini/PE.scala 119:30 123:16 129:16]
  assign io_out_c = {{12{_GEN_7[7]}},_GEN_7}; // @[src/main/scala/gemmini/PE.scala 102:95]
  assign io_out_control_dataflow = io_in_control_dataflow; // @[src/main/scala/gemmini/PE.scala 80:27]
  assign io_out_control_propagate = io_in_control_propagate; // @[src/main/scala/gemmini/PE.scala 81:28]
  assign io_out_control_shift = io_in_control_shift; // @[src/main/scala/gemmini/PE.scala 82:24]
  assign io_out_id = io_in_id; // @[src/main/scala/gemmini/PE.scala 83:13]
  assign io_out_last = io_in_last; // @[src/main/scala/gemmini/PE.scala 84:15]
  assign io_out_valid = io_in_valid; // @[src/main/scala/gemmini/PE.scala 85:16]
  assign mac_unit_io_in_a = io_in_a; // @[src/main/scala/gemmini/PE.scala 87:20]
  assign mac_unit_io_in_b = io_in_control_propagate ? $signed(c2) : $signed(c1); // @[src/main/scala/gemmini/PE.scala 119:30 121:24 127:24]
  assign mac_unit_io_in_c = io_in_b; // @[src/main/scala/gemmini/PE.scala 102:95]
  always @(posedge clock) begin
    c1 <= _GEN_27[7:0];
    c2 <= _GEN_28[7:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c1 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  c2 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_2(
  input         clock,
  input  [7:0]  io_in_a, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [19:0] io_in_b, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [19:0] io_in_d, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [7:0]  io_out_a, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [19:0] io_out_b, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [19:0] io_out_c, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_control_dataflow, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_control_propagate, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [4:0]  io_in_control_shift, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_control_dataflow, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_control_propagate, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [4:0]  io_out_control_shift, // @[src/main/scala/gemmini/PE.scala 35:14]
  input  [1:0]  io_in_id, // @[src/main/scala/gemmini/PE.scala 35:14]
  output [1:0]  io_out_id, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_last, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_last, // @[src/main/scala/gemmini/PE.scala 35:14]
  input         io_in_valid, // @[src/main/scala/gemmini/PE.scala 35:14]
  output        io_out_valid // @[src/main/scala/gemmini/PE.scala 35:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] mac_unit_io_in_a; // @[src/main/scala/gemmini/PE.scala 64:24]
  wire [7:0] mac_unit_io_in_b; // @[src/main/scala/gemmini/PE.scala 64:24]
  wire [19:0] mac_unit_io_in_c; // @[src/main/scala/gemmini/PE.scala 64:24]
  wire [19:0] mac_unit_io_out_d; // @[src/main/scala/gemmini/PE.scala 64:24]
  reg [7:0] c1; // @[src/main/scala/gemmini/PE.scala 70:15]
  reg [7:0] c2; // @[src/main/scala/gemmini/PE.scala 71:15]
  wire [7:0] _GEN_7 = io_in_control_propagate ? $signed(c1) : $signed(c2); // @[src/main/scala/gemmini/PE.scala 119:30 120:16 126:16]
  wire [19:0] _GEN_11 = io_in_control_propagate ? $signed(io_in_d) : $signed({{12{c1[7]}},c1}); // @[src/main/scala/gemmini/PE.scala 119:30 124:10 70:15]
  wire [19:0] _GEN_12 = io_in_control_propagate ? $signed({{12{c2[7]}},c2}) : $signed(io_in_d); // @[src/main/scala/gemmini/PE.scala 119:30 130:10 71:15]
  wire [19:0] _GEN_27 = ~io_in_valid ? $signed({{12{c1[7]}},c1}) : $signed(_GEN_11); // @[src/main/scala/gemmini/PE.scala 141:17 142:8]
  wire [19:0] _GEN_28 = ~io_in_valid ? $signed({{12{c2[7]}},c2}) : $signed(_GEN_12); // @[src/main/scala/gemmini/PE.scala 141:17 143:8]
  MacUnit mac_unit ( // @[src/main/scala/gemmini/PE.scala 64:24]
    .io_in_a(mac_unit_io_in_a),
    .io_in_b(mac_unit_io_in_b),
    .io_in_c(mac_unit_io_in_c),
    .io_out_d(mac_unit_io_out_d)
  );
  assign io_out_a = io_in_a; // @[src/main/scala/gemmini/PE.scala 79:12]
  assign io_out_b = mac_unit_io_out_d; // @[src/main/scala/gemmini/PE.scala 119:30 123:16 129:16]
  assign io_out_c = {{12{_GEN_7[7]}},_GEN_7}; // @[src/main/scala/gemmini/PE.scala 102:95]
  assign io_out_control_dataflow = io_in_control_dataflow; // @[src/main/scala/gemmini/PE.scala 80:27]
  assign io_out_control_propagate = io_in_control_propagate; // @[src/main/scala/gemmini/PE.scala 81:28]
  assign io_out_control_shift = io_in_control_shift; // @[src/main/scala/gemmini/PE.scala 82:24]
  assign io_out_id = io_in_id; // @[src/main/scala/gemmini/PE.scala 83:13]
  assign io_out_last = io_in_last; // @[src/main/scala/gemmini/PE.scala 84:15]
  assign io_out_valid = io_in_valid; // @[src/main/scala/gemmini/PE.scala 85:16]
  assign mac_unit_io_in_a = io_in_a; // @[src/main/scala/gemmini/PE.scala 87:20]
  assign mac_unit_io_in_b = io_in_control_propagate ? $signed(c2) : $signed(c1); // @[src/main/scala/gemmini/PE.scala 119:30 121:24 127:24]
  assign mac_unit_io_in_c = io_in_b; // @[src/main/scala/gemmini/PE.scala 102:95]
  always @(posedge clock) begin
    c1 <= _GEN_27[7:0];
    c2 <= _GEN_28[7:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c1 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  c2 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Tile(
  input         clock,
  input  [7:0]  io_in_a_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [7:0]  io_in_a_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_b_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_b_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_d_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_d_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_0_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_0_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [4:0]  io_in_control_0_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_1_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_1_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [4:0]  io_in_control_1_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [1:0]  io_in_id_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [1:0]  io_in_id_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_last_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_last_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [7:0]  io_out_a_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [7:0]  io_out_a_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_c_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_c_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_b_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_b_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_0_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_0_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [4:0]  io_out_control_0_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_1_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_1_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [4:0]  io_out_control_1_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [1:0]  io_out_id_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [1:0]  io_out_id_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_last_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_last_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_valid_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_valid_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_valid_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_valid_1 // @[src/main/scala/gemmini/Tile.scala 17:14]
);
  wire  tile_0_0_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_0_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_0_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_0_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_1_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_1_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_1_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_0_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_0_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_0_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_1_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_1_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_1_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  PE tile_0_0 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_0_0_clock),
    .io_in_a(tile_0_0_io_in_a),
    .io_in_b(tile_0_0_io_in_b),
    .io_in_d(tile_0_0_io_in_d),
    .io_out_a(tile_0_0_io_out_a),
    .io_out_b(tile_0_0_io_out_b),
    .io_out_c(tile_0_0_io_out_c),
    .io_in_control_dataflow(tile_0_0_io_in_control_dataflow),
    .io_in_control_propagate(tile_0_0_io_in_control_propagate),
    .io_in_control_shift(tile_0_0_io_in_control_shift),
    .io_out_control_dataflow(tile_0_0_io_out_control_dataflow),
    .io_out_control_propagate(tile_0_0_io_out_control_propagate),
    .io_out_control_shift(tile_0_0_io_out_control_shift),
    .io_in_id(tile_0_0_io_in_id),
    .io_out_id(tile_0_0_io_out_id),
    .io_in_last(tile_0_0_io_in_last),
    .io_out_last(tile_0_0_io_out_last),
    .io_in_valid(tile_0_0_io_in_valid),
    .io_out_valid(tile_0_0_io_out_valid)
  );
  PE tile_0_1 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_0_1_clock),
    .io_in_a(tile_0_1_io_in_a),
    .io_in_b(tile_0_1_io_in_b),
    .io_in_d(tile_0_1_io_in_d),
    .io_out_a(tile_0_1_io_out_a),
    .io_out_b(tile_0_1_io_out_b),
    .io_out_c(tile_0_1_io_out_c),
    .io_in_control_dataflow(tile_0_1_io_in_control_dataflow),
    .io_in_control_propagate(tile_0_1_io_in_control_propagate),
    .io_in_control_shift(tile_0_1_io_in_control_shift),
    .io_out_control_dataflow(tile_0_1_io_out_control_dataflow),
    .io_out_control_propagate(tile_0_1_io_out_control_propagate),
    .io_out_control_shift(tile_0_1_io_out_control_shift),
    .io_in_id(tile_0_1_io_in_id),
    .io_out_id(tile_0_1_io_out_id),
    .io_in_last(tile_0_1_io_in_last),
    .io_out_last(tile_0_1_io_out_last),
    .io_in_valid(tile_0_1_io_in_valid),
    .io_out_valid(tile_0_1_io_out_valid)
  );
  PE_2 tile_1_0 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_1_0_clock),
    .io_in_a(tile_1_0_io_in_a),
    .io_in_b(tile_1_0_io_in_b),
    .io_in_d(tile_1_0_io_in_d),
    .io_out_a(tile_1_0_io_out_a),
    .io_out_b(tile_1_0_io_out_b),
    .io_out_c(tile_1_0_io_out_c),
    .io_in_control_dataflow(tile_1_0_io_in_control_dataflow),
    .io_in_control_propagate(tile_1_0_io_in_control_propagate),
    .io_in_control_shift(tile_1_0_io_in_control_shift),
    .io_out_control_dataflow(tile_1_0_io_out_control_dataflow),
    .io_out_control_propagate(tile_1_0_io_out_control_propagate),
    .io_out_control_shift(tile_1_0_io_out_control_shift),
    .io_in_id(tile_1_0_io_in_id),
    .io_out_id(tile_1_0_io_out_id),
    .io_in_last(tile_1_0_io_in_last),
    .io_out_last(tile_1_0_io_out_last),
    .io_in_valid(tile_1_0_io_in_valid),
    .io_out_valid(tile_1_0_io_out_valid)
  );
  PE_2 tile_1_1 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_1_1_clock),
    .io_in_a(tile_1_1_io_in_a),
    .io_in_b(tile_1_1_io_in_b),
    .io_in_d(tile_1_1_io_in_d),
    .io_out_a(tile_1_1_io_out_a),
    .io_out_b(tile_1_1_io_out_b),
    .io_out_c(tile_1_1_io_out_c),
    .io_in_control_dataflow(tile_1_1_io_in_control_dataflow),
    .io_in_control_propagate(tile_1_1_io_in_control_propagate),
    .io_in_control_shift(tile_1_1_io_in_control_shift),
    .io_out_control_dataflow(tile_1_1_io_out_control_dataflow),
    .io_out_control_propagate(tile_1_1_io_out_control_propagate),
    .io_out_control_shift(tile_1_1_io_out_control_shift),
    .io_in_id(tile_1_1_io_in_id),
    .io_out_id(tile_1_1_io_out_id),
    .io_in_last(tile_1_1_io_in_last),
    .io_out_last(tile_1_1_io_out_last),
    .io_in_valid(tile_1_1_io_in_valid),
    .io_out_valid(tile_1_1_io_out_valid)
  );
  assign io_out_a_0 = tile_0_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 130:17]
  assign io_out_a_1 = tile_1_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 130:17]
  assign io_out_c_0 = tile_1_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 111:17]
  assign io_out_c_1 = tile_1_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 111:17]
  assign io_out_b_0 = tile_1_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 117:17]
  assign io_out_b_1 = tile_1_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 117:17]
  assign io_out_control_0_dataflow = tile_1_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_0_propagate = tile_1_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_0_shift = tile_1_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_1_dataflow = tile_1_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_1_propagate = tile_1_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_1_shift = tile_1_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_id_0 = tile_1_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 113:18]
  assign io_out_id_1 = tile_1_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 113:18]
  assign io_out_last_0 = tile_1_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 114:20]
  assign io_out_last_1 = tile_1_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 114:20]
  assign io_out_valid_0 = tile_1_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 115:21]
  assign io_out_valid_1 = tile_1_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 115:21]
  assign tile_0_0_clock = clock;
  assign tile_0_0_io_in_a = io_in_a_0; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_0_0_io_in_b = io_in_b_0; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_0_0_io_in_d = io_in_d_0; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_0_0_io_in_control_dataflow = io_in_control_0_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_0_io_in_control_propagate = io_in_control_0_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_0_io_in_control_shift = io_in_control_0_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_0_io_in_id = io_in_id_0; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_0_0_io_in_last = io_in_last_0; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_0_0_io_in_valid = io_in_valid_0; // @[src/main/scala/gemmini/Tile.scala 86:24]
  assign tile_0_1_clock = clock;
  assign tile_0_1_io_in_a = tile_0_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_0_1_io_in_b = io_in_b_1; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_0_1_io_in_d = io_in_d_1; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_0_1_io_in_control_dataflow = io_in_control_1_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_1_io_in_control_propagate = io_in_control_1_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_1_io_in_control_shift = io_in_control_1_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_1_io_in_id = io_in_id_1; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_0_1_io_in_last = io_in_last_1; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_0_1_io_in_valid = io_in_valid_1; // @[src/main/scala/gemmini/Tile.scala 86:24]
  assign tile_1_0_clock = clock;
  assign tile_1_0_io_in_a = io_in_a_1; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_1_0_io_in_b = tile_0_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_1_0_io_in_d = tile_0_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_1_0_io_in_control_dataflow = tile_0_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_0_io_in_control_propagate = tile_0_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_0_io_in_control_shift = tile_0_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_0_io_in_id = tile_0_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_1_0_io_in_last = tile_0_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_1_0_io_in_valid = tile_0_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 86:24]
  assign tile_1_1_clock = clock;
  assign tile_1_1_io_in_a = tile_1_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_1_1_io_in_b = tile_0_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_1_1_io_in_d = tile_0_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_1_1_io_in_control_dataflow = tile_0_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_1_io_in_control_propagate = tile_0_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_1_io_in_control_shift = tile_0_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_1_io_in_id = tile_0_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_1_1_io_in_last = tile_0_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_1_1_io_in_valid = tile_0_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 86:24]
endmodule
module Tile_240(
  input         clock,
  input  [7:0]  io_in_a_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [7:0]  io_in_a_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_b_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_b_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_d_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [19:0] io_in_d_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_0_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_0_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [4:0]  io_in_control_0_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_1_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_control_1_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [4:0]  io_in_control_1_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [1:0]  io_in_id_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input  [1:0]  io_in_id_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_last_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_last_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [7:0]  io_out_a_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [7:0]  io_out_a_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_c_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_c_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_b_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [19:0] io_out_b_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_0_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_0_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [4:0]  io_out_control_0_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_1_dataflow, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_control_1_propagate, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [4:0]  io_out_control_1_shift, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [1:0]  io_out_id_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output [1:0]  io_out_id_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_last_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_last_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_valid_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  input         io_in_valid_1, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_valid_0, // @[src/main/scala/gemmini/Tile.scala 17:14]
  output        io_out_valid_1 // @[src/main/scala/gemmini/Tile.scala 17:14]
);
  wire  tile_0_0_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_0_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_0_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_0_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_1_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_0_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_0_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_1_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_0_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_1_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_0_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_0_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_0_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_0_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_0_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_clock; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_1_io_in_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_in_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_in_d; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [7:0] tile_1_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [19:0] tile_1_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_1_io_in_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [4:0] tile_1_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_1_io_in_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire [1:0] tile_1_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_in_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  wire  tile_1_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 42:44]
  PE tile_0_0 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_0_0_clock),
    .io_in_a(tile_0_0_io_in_a),
    .io_in_b(tile_0_0_io_in_b),
    .io_in_d(tile_0_0_io_in_d),
    .io_out_a(tile_0_0_io_out_a),
    .io_out_b(tile_0_0_io_out_b),
    .io_out_c(tile_0_0_io_out_c),
    .io_in_control_dataflow(tile_0_0_io_in_control_dataflow),
    .io_in_control_propagate(tile_0_0_io_in_control_propagate),
    .io_in_control_shift(tile_0_0_io_in_control_shift),
    .io_out_control_dataflow(tile_0_0_io_out_control_dataflow),
    .io_out_control_propagate(tile_0_0_io_out_control_propagate),
    .io_out_control_shift(tile_0_0_io_out_control_shift),
    .io_in_id(tile_0_0_io_in_id),
    .io_out_id(tile_0_0_io_out_id),
    .io_in_last(tile_0_0_io_in_last),
    .io_out_last(tile_0_0_io_out_last),
    .io_in_valid(tile_0_0_io_in_valid),
    .io_out_valid(tile_0_0_io_out_valid)
  );
  PE tile_0_1 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_0_1_clock),
    .io_in_a(tile_0_1_io_in_a),
    .io_in_b(tile_0_1_io_in_b),
    .io_in_d(tile_0_1_io_in_d),
    .io_out_a(tile_0_1_io_out_a),
    .io_out_b(tile_0_1_io_out_b),
    .io_out_c(tile_0_1_io_out_c),
    .io_in_control_dataflow(tile_0_1_io_in_control_dataflow),
    .io_in_control_propagate(tile_0_1_io_in_control_propagate),
    .io_in_control_shift(tile_0_1_io_in_control_shift),
    .io_out_control_dataflow(tile_0_1_io_out_control_dataflow),
    .io_out_control_propagate(tile_0_1_io_out_control_propagate),
    .io_out_control_shift(tile_0_1_io_out_control_shift),
    .io_in_id(tile_0_1_io_in_id),
    .io_out_id(tile_0_1_io_out_id),
    .io_in_last(tile_0_1_io_in_last),
    .io_out_last(tile_0_1_io_out_last),
    .io_in_valid(tile_0_1_io_in_valid),
    .io_out_valid(tile_0_1_io_out_valid)
  );
  PE_2 tile_1_0 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_1_0_clock),
    .io_in_a(tile_1_0_io_in_a),
    .io_in_b(tile_1_0_io_in_b),
    .io_in_d(tile_1_0_io_in_d),
    .io_out_a(tile_1_0_io_out_a),
    .io_out_b(tile_1_0_io_out_b),
    .io_out_c(tile_1_0_io_out_c),
    .io_in_control_dataflow(tile_1_0_io_in_control_dataflow),
    .io_in_control_propagate(tile_1_0_io_in_control_propagate),
    .io_in_control_shift(tile_1_0_io_in_control_shift),
    .io_out_control_dataflow(tile_1_0_io_out_control_dataflow),
    .io_out_control_propagate(tile_1_0_io_out_control_propagate),
    .io_out_control_shift(tile_1_0_io_out_control_shift),
    .io_in_id(tile_1_0_io_in_id),
    .io_out_id(tile_1_0_io_out_id),
    .io_in_last(tile_1_0_io_in_last),
    .io_out_last(tile_1_0_io_out_last),
    .io_in_valid(tile_1_0_io_in_valid),
    .io_out_valid(tile_1_0_io_out_valid)
  );
  PE_2 tile_1_1 ( // @[src/main/scala/gemmini/Tile.scala 42:44]
    .clock(tile_1_1_clock),
    .io_in_a(tile_1_1_io_in_a),
    .io_in_b(tile_1_1_io_in_b),
    .io_in_d(tile_1_1_io_in_d),
    .io_out_a(tile_1_1_io_out_a),
    .io_out_b(tile_1_1_io_out_b),
    .io_out_c(tile_1_1_io_out_c),
    .io_in_control_dataflow(tile_1_1_io_in_control_dataflow),
    .io_in_control_propagate(tile_1_1_io_in_control_propagate),
    .io_in_control_shift(tile_1_1_io_in_control_shift),
    .io_out_control_dataflow(tile_1_1_io_out_control_dataflow),
    .io_out_control_propagate(tile_1_1_io_out_control_propagate),
    .io_out_control_shift(tile_1_1_io_out_control_shift),
    .io_in_id(tile_1_1_io_in_id),
    .io_out_id(tile_1_1_io_out_id),
    .io_in_last(tile_1_1_io_in_last),
    .io_out_last(tile_1_1_io_out_last),
    .io_in_valid(tile_1_1_io_in_valid),
    .io_out_valid(tile_1_1_io_out_valid)
  );
  assign io_out_a_0 = tile_0_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 130:17]
  assign io_out_a_1 = tile_1_1_io_out_a; // @[src/main/scala/gemmini/Tile.scala 130:17]
  assign io_out_c_0 = tile_1_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 111:17]
  assign io_out_c_1 = tile_1_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 111:17]
  assign io_out_b_0 = tile_1_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 117:17]
  assign io_out_b_1 = tile_1_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 117:17]
  assign io_out_control_0_dataflow = tile_1_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_0_propagate = tile_1_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_0_shift = tile_1_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_1_dataflow = tile_1_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_1_propagate = tile_1_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_control_1_shift = tile_1_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 112:23]
  assign io_out_id_0 = tile_1_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 113:18]
  assign io_out_id_1 = tile_1_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 113:18]
  assign io_out_last_0 = tile_1_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 114:20]
  assign io_out_last_1 = tile_1_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 114:20]
  assign io_out_valid_0 = tile_1_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 115:21]
  assign io_out_valid_1 = tile_1_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 115:21]
  assign tile_0_0_clock = clock;
  assign tile_0_0_io_in_a = io_in_a_0; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_0_0_io_in_b = io_in_b_0; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_0_0_io_in_d = io_in_d_0; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_0_0_io_in_control_dataflow = io_in_control_0_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_0_io_in_control_propagate = io_in_control_0_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_0_io_in_control_shift = io_in_control_0_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_0_io_in_id = io_in_id_0; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_0_0_io_in_last = io_in_last_0; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_0_0_io_in_valid = io_in_valid_0; // @[src/main/scala/gemmini/Tile.scala 86:24]
  assign tile_0_1_clock = clock;
  assign tile_0_1_io_in_a = tile_0_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_0_1_io_in_b = io_in_b_1; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_0_1_io_in_d = io_in_d_1; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_0_1_io_in_control_dataflow = io_in_control_1_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_1_io_in_control_propagate = io_in_control_1_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_1_io_in_control_shift = io_in_control_1_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_0_1_io_in_id = io_in_id_1; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_0_1_io_in_last = io_in_last_1; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_0_1_io_in_valid = io_in_valid_1; // @[src/main/scala/gemmini/Tile.scala 86:24]
  assign tile_1_0_clock = clock;
  assign tile_1_0_io_in_a = io_in_a_1; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_1_0_io_in_b = tile_0_0_io_out_b; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_1_0_io_in_d = tile_0_0_io_out_c; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_1_0_io_in_control_dataflow = tile_0_0_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_0_io_in_control_propagate = tile_0_0_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_0_io_in_control_shift = tile_0_0_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_0_io_in_id = tile_0_0_io_out_id; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_1_0_io_in_last = tile_0_0_io_out_last; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_1_0_io_in_valid = tile_0_0_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 86:24]
  assign tile_1_1_clock = clock;
  assign tile_1_1_io_in_a = tile_1_0_io_out_a; // @[src/main/scala/gemmini/Tile.scala 50:20]
  assign tile_1_1_io_in_b = tile_0_1_io_out_b; // @[src/main/scala/gemmini/Tile.scala 59:20]
  assign tile_1_1_io_in_d = tile_0_1_io_out_c; // @[src/main/scala/gemmini/Tile.scala 68:20]
  assign tile_1_1_io_in_control_dataflow = tile_0_1_io_out_control_dataflow; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_1_io_in_control_propagate = tile_0_1_io_out_control_propagate; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_1_io_in_control_shift = tile_0_1_io_out_control_shift; // @[src/main/scala/gemmini/Tile.scala 77:26]
  assign tile_1_1_io_in_id = tile_0_1_io_out_id; // @[src/main/scala/gemmini/Tile.scala 95:21]
  assign tile_1_1_io_in_last = tile_0_1_io_out_last; // @[src/main/scala/gemmini/Tile.scala 104:23]
  assign tile_1_1_io_in_valid = tile_0_1_io_out_valid; // @[src/main/scala/gemmini/Tile.scala 86:24]
endmodule
module Mesh(
  input         clock,
  input  [7:0]  io_in_a_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_a_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_b_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [7:0]  io_in_d_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_0_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_0_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_0_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_0_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_0_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_0_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_1_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_1_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_1_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_1_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_1_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_1_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_2_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_2_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_2_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_2_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_2_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_2_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_3_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_3_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_3_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_3_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_3_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_3_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_4_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_4_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_4_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_4_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_4_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_4_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_5_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_5_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_5_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_5_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_5_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_5_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_6_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_6_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_6_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_6_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_6_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_6_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_7_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_7_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_7_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_7_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_7_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_7_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_8_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_8_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_8_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_8_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_8_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_8_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_9_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_9_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_9_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_9_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_9_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_9_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_10_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_10_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_10_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_10_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_10_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_10_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_11_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_11_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_11_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_11_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_11_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_11_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_12_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_12_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_12_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_12_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_12_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_12_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_13_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_13_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_13_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_13_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_13_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_13_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_14_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_14_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_14_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_14_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_14_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_14_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_15_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_15_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_15_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_15_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_control_15_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [4:0]  io_in_control_15_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input  [1:0]  io_in_id_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_last_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_b_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [19:0] io_out_c_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  input         io_in_valid_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_valid_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_0_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_0_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_0_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_0_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_0_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_0_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_1_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_1_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_1_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_1_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_1_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_1_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_2_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_2_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_2_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_2_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_2_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_2_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_3_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_3_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_3_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_3_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_3_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_3_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_4_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_4_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_4_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_4_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_4_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_4_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_5_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_5_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_5_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_5_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_5_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_5_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_6_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_6_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_6_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_6_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_6_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_6_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_7_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_7_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_7_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_7_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_7_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_7_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_8_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_8_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_8_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_8_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_8_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_8_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_9_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_9_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_9_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_9_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_9_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_9_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_10_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_10_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_10_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_10_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_10_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_10_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_11_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_11_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_11_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_11_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_11_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_11_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_12_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_12_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_12_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_12_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_12_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_12_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_13_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_13_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_13_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_13_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_13_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_13_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_14_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_14_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_14_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_14_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_14_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_14_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_15_0_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_15_0_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_15_0_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_15_1_dataflow, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_control_15_1_propagate, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [4:0]  io_out_control_15_1_shift, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output [1:0]  io_out_id_15_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_0_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_0_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_1_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_1_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_2_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_2_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_3_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_3_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_4_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_4_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_5_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_5_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_6_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_6_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_7_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_7_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_8_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_8_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_9_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_9_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_10_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_10_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_11_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_11_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_12_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_12_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_13_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_13_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_14_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_14_1, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_15_0, // @[src/main/scala/gemmini/Mesh.scala 22:14]
  output        io_out_last_15_1 // @[src/main/scala/gemmini/Mesh.scala 22:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [31:0] _RAND_2817;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
  reg [31:0] _RAND_2841;
  reg [31:0] _RAND_2842;
  reg [31:0] _RAND_2843;
  reg [31:0] _RAND_2844;
  reg [31:0] _RAND_2845;
  reg [31:0] _RAND_2846;
  reg [31:0] _RAND_2847;
  reg [31:0] _RAND_2848;
  reg [31:0] _RAND_2849;
  reg [31:0] _RAND_2850;
  reg [31:0] _RAND_2851;
  reg [31:0] _RAND_2852;
  reg [31:0] _RAND_2853;
  reg [31:0] _RAND_2854;
  reg [31:0] _RAND_2855;
  reg [31:0] _RAND_2856;
  reg [31:0] _RAND_2857;
  reg [31:0] _RAND_2858;
  reg [31:0] _RAND_2859;
  reg [31:0] _RAND_2860;
  reg [31:0] _RAND_2861;
  reg [31:0] _RAND_2862;
  reg [31:0] _RAND_2863;
  reg [31:0] _RAND_2864;
  reg [31:0] _RAND_2865;
  reg [31:0] _RAND_2866;
  reg [31:0] _RAND_2867;
  reg [31:0] _RAND_2868;
  reg [31:0] _RAND_2869;
  reg [31:0] _RAND_2870;
  reg [31:0] _RAND_2871;
  reg [31:0] _RAND_2872;
  reg [31:0] _RAND_2873;
  reg [31:0] _RAND_2874;
  reg [31:0] _RAND_2875;
  reg [31:0] _RAND_2876;
  reg [31:0] _RAND_2877;
  reg [31:0] _RAND_2878;
  reg [31:0] _RAND_2879;
  reg [31:0] _RAND_2880;
  reg [31:0] _RAND_2881;
  reg [31:0] _RAND_2882;
  reg [31:0] _RAND_2883;
  reg [31:0] _RAND_2884;
  reg [31:0] _RAND_2885;
  reg [31:0] _RAND_2886;
  reg [31:0] _RAND_2887;
  reg [31:0] _RAND_2888;
  reg [31:0] _RAND_2889;
  reg [31:0] _RAND_2890;
  reg [31:0] _RAND_2891;
  reg [31:0] _RAND_2892;
  reg [31:0] _RAND_2893;
  reg [31:0] _RAND_2894;
  reg [31:0] _RAND_2895;
  reg [31:0] _RAND_2896;
  reg [31:0] _RAND_2897;
  reg [31:0] _RAND_2898;
  reg [31:0] _RAND_2899;
  reg [31:0] _RAND_2900;
  reg [31:0] _RAND_2901;
  reg [31:0] _RAND_2902;
  reg [31:0] _RAND_2903;
  reg [31:0] _RAND_2904;
  reg [31:0] _RAND_2905;
  reg [31:0] _RAND_2906;
  reg [31:0] _RAND_2907;
  reg [31:0] _RAND_2908;
  reg [31:0] _RAND_2909;
  reg [31:0] _RAND_2910;
  reg [31:0] _RAND_2911;
  reg [31:0] _RAND_2912;
  reg [31:0] _RAND_2913;
  reg [31:0] _RAND_2914;
  reg [31:0] _RAND_2915;
  reg [31:0] _RAND_2916;
  reg [31:0] _RAND_2917;
  reg [31:0] _RAND_2918;
  reg [31:0] _RAND_2919;
  reg [31:0] _RAND_2920;
  reg [31:0] _RAND_2921;
  reg [31:0] _RAND_2922;
  reg [31:0] _RAND_2923;
  reg [31:0] _RAND_2924;
  reg [31:0] _RAND_2925;
  reg [31:0] _RAND_2926;
  reg [31:0] _RAND_2927;
  reg [31:0] _RAND_2928;
  reg [31:0] _RAND_2929;
  reg [31:0] _RAND_2930;
  reg [31:0] _RAND_2931;
  reg [31:0] _RAND_2932;
  reg [31:0] _RAND_2933;
  reg [31:0] _RAND_2934;
  reg [31:0] _RAND_2935;
  reg [31:0] _RAND_2936;
  reg [31:0] _RAND_2937;
  reg [31:0] _RAND_2938;
  reg [31:0] _RAND_2939;
  reg [31:0] _RAND_2940;
  reg [31:0] _RAND_2941;
  reg [31:0] _RAND_2942;
  reg [31:0] _RAND_2943;
  reg [31:0] _RAND_2944;
  reg [31:0] _RAND_2945;
  reg [31:0] _RAND_2946;
  reg [31:0] _RAND_2947;
  reg [31:0] _RAND_2948;
  reg [31:0] _RAND_2949;
  reg [31:0] _RAND_2950;
  reg [31:0] _RAND_2951;
  reg [31:0] _RAND_2952;
  reg [31:0] _RAND_2953;
  reg [31:0] _RAND_2954;
  reg [31:0] _RAND_2955;
  reg [31:0] _RAND_2956;
  reg [31:0] _RAND_2957;
  reg [31:0] _RAND_2958;
  reg [31:0] _RAND_2959;
  reg [31:0] _RAND_2960;
  reg [31:0] _RAND_2961;
  reg [31:0] _RAND_2962;
  reg [31:0] _RAND_2963;
  reg [31:0] _RAND_2964;
  reg [31:0] _RAND_2965;
  reg [31:0] _RAND_2966;
  reg [31:0] _RAND_2967;
  reg [31:0] _RAND_2968;
  reg [31:0] _RAND_2969;
  reg [31:0] _RAND_2970;
  reg [31:0] _RAND_2971;
  reg [31:0] _RAND_2972;
  reg [31:0] _RAND_2973;
  reg [31:0] _RAND_2974;
  reg [31:0] _RAND_2975;
  reg [31:0] _RAND_2976;
  reg [31:0] _RAND_2977;
  reg [31:0] _RAND_2978;
  reg [31:0] _RAND_2979;
  reg [31:0] _RAND_2980;
  reg [31:0] _RAND_2981;
  reg [31:0] _RAND_2982;
  reg [31:0] _RAND_2983;
  reg [31:0] _RAND_2984;
  reg [31:0] _RAND_2985;
  reg [31:0] _RAND_2986;
  reg [31:0] _RAND_2987;
  reg [31:0] _RAND_2988;
  reg [31:0] _RAND_2989;
  reg [31:0] _RAND_2990;
  reg [31:0] _RAND_2991;
  reg [31:0] _RAND_2992;
  reg [31:0] _RAND_2993;
  reg [31:0] _RAND_2994;
  reg [31:0] _RAND_2995;
  reg [31:0] _RAND_2996;
  reg [31:0] _RAND_2997;
  reg [31:0] _RAND_2998;
  reg [31:0] _RAND_2999;
  reg [31:0] _RAND_3000;
  reg [31:0] _RAND_3001;
  reg [31:0] _RAND_3002;
  reg [31:0] _RAND_3003;
  reg [31:0] _RAND_3004;
  reg [31:0] _RAND_3005;
  reg [31:0] _RAND_3006;
  reg [31:0] _RAND_3007;
  reg [31:0] _RAND_3008;
  reg [31:0] _RAND_3009;
  reg [31:0] _RAND_3010;
  reg [31:0] _RAND_3011;
  reg [31:0] _RAND_3012;
  reg [31:0] _RAND_3013;
  reg [31:0] _RAND_3014;
  reg [31:0] _RAND_3015;
  reg [31:0] _RAND_3016;
  reg [31:0] _RAND_3017;
  reg [31:0] _RAND_3018;
  reg [31:0] _RAND_3019;
  reg [31:0] _RAND_3020;
  reg [31:0] _RAND_3021;
  reg [31:0] _RAND_3022;
  reg [31:0] _RAND_3023;
  reg [31:0] _RAND_3024;
  reg [31:0] _RAND_3025;
  reg [31:0] _RAND_3026;
  reg [31:0] _RAND_3027;
  reg [31:0] _RAND_3028;
  reg [31:0] _RAND_3029;
  reg [31:0] _RAND_3030;
  reg [31:0] _RAND_3031;
  reg [31:0] _RAND_3032;
  reg [31:0] _RAND_3033;
  reg [31:0] _RAND_3034;
  reg [31:0] _RAND_3035;
  reg [31:0] _RAND_3036;
  reg [31:0] _RAND_3037;
  reg [31:0] _RAND_3038;
  reg [31:0] _RAND_3039;
  reg [31:0] _RAND_3040;
  reg [31:0] _RAND_3041;
  reg [31:0] _RAND_3042;
  reg [31:0] _RAND_3043;
  reg [31:0] _RAND_3044;
  reg [31:0] _RAND_3045;
  reg [31:0] _RAND_3046;
  reg [31:0] _RAND_3047;
  reg [31:0] _RAND_3048;
  reg [31:0] _RAND_3049;
  reg [31:0] _RAND_3050;
  reg [31:0] _RAND_3051;
  reg [31:0] _RAND_3052;
  reg [31:0] _RAND_3053;
  reg [31:0] _RAND_3054;
  reg [31:0] _RAND_3055;
  reg [31:0] _RAND_3056;
  reg [31:0] _RAND_3057;
  reg [31:0] _RAND_3058;
  reg [31:0] _RAND_3059;
  reg [31:0] _RAND_3060;
  reg [31:0] _RAND_3061;
  reg [31:0] _RAND_3062;
  reg [31:0] _RAND_3063;
  reg [31:0] _RAND_3064;
  reg [31:0] _RAND_3065;
  reg [31:0] _RAND_3066;
  reg [31:0] _RAND_3067;
  reg [31:0] _RAND_3068;
  reg [31:0] _RAND_3069;
  reg [31:0] _RAND_3070;
  reg [31:0] _RAND_3071;
  reg [31:0] _RAND_3072;
  reg [31:0] _RAND_3073;
  reg [31:0] _RAND_3074;
  reg [31:0] _RAND_3075;
  reg [31:0] _RAND_3076;
  reg [31:0] _RAND_3077;
  reg [31:0] _RAND_3078;
  reg [31:0] _RAND_3079;
  reg [31:0] _RAND_3080;
  reg [31:0] _RAND_3081;
  reg [31:0] _RAND_3082;
  reg [31:0] _RAND_3083;
  reg [31:0] _RAND_3084;
  reg [31:0] _RAND_3085;
  reg [31:0] _RAND_3086;
  reg [31:0] _RAND_3087;
  reg [31:0] _RAND_3088;
  reg [31:0] _RAND_3089;
  reg [31:0] _RAND_3090;
  reg [31:0] _RAND_3091;
  reg [31:0] _RAND_3092;
  reg [31:0] _RAND_3093;
  reg [31:0] _RAND_3094;
  reg [31:0] _RAND_3095;
  reg [31:0] _RAND_3096;
  reg [31:0] _RAND_3097;
  reg [31:0] _RAND_3098;
  reg [31:0] _RAND_3099;
  reg [31:0] _RAND_3100;
  reg [31:0] _RAND_3101;
  reg [31:0] _RAND_3102;
  reg [31:0] _RAND_3103;
  reg [31:0] _RAND_3104;
  reg [31:0] _RAND_3105;
  reg [31:0] _RAND_3106;
  reg [31:0] _RAND_3107;
  reg [31:0] _RAND_3108;
  reg [31:0] _RAND_3109;
  reg [31:0] _RAND_3110;
  reg [31:0] _RAND_3111;
  reg [31:0] _RAND_3112;
  reg [31:0] _RAND_3113;
  reg [31:0] _RAND_3114;
  reg [31:0] _RAND_3115;
  reg [31:0] _RAND_3116;
  reg [31:0] _RAND_3117;
  reg [31:0] _RAND_3118;
  reg [31:0] _RAND_3119;
  reg [31:0] _RAND_3120;
  reg [31:0] _RAND_3121;
  reg [31:0] _RAND_3122;
  reg [31:0] _RAND_3123;
  reg [31:0] _RAND_3124;
  reg [31:0] _RAND_3125;
  reg [31:0] _RAND_3126;
  reg [31:0] _RAND_3127;
  reg [31:0] _RAND_3128;
  reg [31:0] _RAND_3129;
  reg [31:0] _RAND_3130;
  reg [31:0] _RAND_3131;
  reg [31:0] _RAND_3132;
  reg [31:0] _RAND_3133;
  reg [31:0] _RAND_3134;
  reg [31:0] _RAND_3135;
  reg [31:0] _RAND_3136;
  reg [31:0] _RAND_3137;
  reg [31:0] _RAND_3138;
  reg [31:0] _RAND_3139;
  reg [31:0] _RAND_3140;
  reg [31:0] _RAND_3141;
  reg [31:0] _RAND_3142;
  reg [31:0] _RAND_3143;
  reg [31:0] _RAND_3144;
  reg [31:0] _RAND_3145;
  reg [31:0] _RAND_3146;
  reg [31:0] _RAND_3147;
  reg [31:0] _RAND_3148;
  reg [31:0] _RAND_3149;
  reg [31:0] _RAND_3150;
  reg [31:0] _RAND_3151;
  reg [31:0] _RAND_3152;
  reg [31:0] _RAND_3153;
  reg [31:0] _RAND_3154;
  reg [31:0] _RAND_3155;
  reg [31:0] _RAND_3156;
  reg [31:0] _RAND_3157;
  reg [31:0] _RAND_3158;
  reg [31:0] _RAND_3159;
  reg [31:0] _RAND_3160;
  reg [31:0] _RAND_3161;
  reg [31:0] _RAND_3162;
  reg [31:0] _RAND_3163;
  reg [31:0] _RAND_3164;
  reg [31:0] _RAND_3165;
  reg [31:0] _RAND_3166;
  reg [31:0] _RAND_3167;
  reg [31:0] _RAND_3168;
  reg [31:0] _RAND_3169;
  reg [31:0] _RAND_3170;
  reg [31:0] _RAND_3171;
  reg [31:0] _RAND_3172;
  reg [31:0] _RAND_3173;
  reg [31:0] _RAND_3174;
  reg [31:0] _RAND_3175;
  reg [31:0] _RAND_3176;
  reg [31:0] _RAND_3177;
  reg [31:0] _RAND_3178;
  reg [31:0] _RAND_3179;
  reg [31:0] _RAND_3180;
  reg [31:0] _RAND_3181;
  reg [31:0] _RAND_3182;
  reg [31:0] _RAND_3183;
  reg [31:0] _RAND_3184;
  reg [31:0] _RAND_3185;
  reg [31:0] _RAND_3186;
  reg [31:0] _RAND_3187;
  reg [31:0] _RAND_3188;
  reg [31:0] _RAND_3189;
  reg [31:0] _RAND_3190;
  reg [31:0] _RAND_3191;
  reg [31:0] _RAND_3192;
  reg [31:0] _RAND_3193;
  reg [31:0] _RAND_3194;
  reg [31:0] _RAND_3195;
  reg [31:0] _RAND_3196;
  reg [31:0] _RAND_3197;
  reg [31:0] _RAND_3198;
  reg [31:0] _RAND_3199;
  reg [31:0] _RAND_3200;
  reg [31:0] _RAND_3201;
  reg [31:0] _RAND_3202;
  reg [31:0] _RAND_3203;
  reg [31:0] _RAND_3204;
  reg [31:0] _RAND_3205;
  reg [31:0] _RAND_3206;
  reg [31:0] _RAND_3207;
  reg [31:0] _RAND_3208;
  reg [31:0] _RAND_3209;
  reg [31:0] _RAND_3210;
  reg [31:0] _RAND_3211;
  reg [31:0] _RAND_3212;
  reg [31:0] _RAND_3213;
  reg [31:0] _RAND_3214;
  reg [31:0] _RAND_3215;
  reg [31:0] _RAND_3216;
  reg [31:0] _RAND_3217;
  reg [31:0] _RAND_3218;
  reg [31:0] _RAND_3219;
  reg [31:0] _RAND_3220;
  reg [31:0] _RAND_3221;
  reg [31:0] _RAND_3222;
  reg [31:0] _RAND_3223;
  reg [31:0] _RAND_3224;
  reg [31:0] _RAND_3225;
  reg [31:0] _RAND_3226;
  reg [31:0] _RAND_3227;
  reg [31:0] _RAND_3228;
  reg [31:0] _RAND_3229;
  reg [31:0] _RAND_3230;
  reg [31:0] _RAND_3231;
  reg [31:0] _RAND_3232;
  reg [31:0] _RAND_3233;
  reg [31:0] _RAND_3234;
  reg [31:0] _RAND_3235;
  reg [31:0] _RAND_3236;
  reg [31:0] _RAND_3237;
  reg [31:0] _RAND_3238;
  reg [31:0] _RAND_3239;
  reg [31:0] _RAND_3240;
  reg [31:0] _RAND_3241;
  reg [31:0] _RAND_3242;
  reg [31:0] _RAND_3243;
  reg [31:0] _RAND_3244;
  reg [31:0] _RAND_3245;
  reg [31:0] _RAND_3246;
  reg [31:0] _RAND_3247;
  reg [31:0] _RAND_3248;
  reg [31:0] _RAND_3249;
  reg [31:0] _RAND_3250;
  reg [31:0] _RAND_3251;
  reg [31:0] _RAND_3252;
  reg [31:0] _RAND_3253;
  reg [31:0] _RAND_3254;
  reg [31:0] _RAND_3255;
  reg [31:0] _RAND_3256;
  reg [31:0] _RAND_3257;
  reg [31:0] _RAND_3258;
  reg [31:0] _RAND_3259;
  reg [31:0] _RAND_3260;
  reg [31:0] _RAND_3261;
  reg [31:0] _RAND_3262;
  reg [31:0] _RAND_3263;
  reg [31:0] _RAND_3264;
  reg [31:0] _RAND_3265;
  reg [31:0] _RAND_3266;
  reg [31:0] _RAND_3267;
  reg [31:0] _RAND_3268;
  reg [31:0] _RAND_3269;
  reg [31:0] _RAND_3270;
  reg [31:0] _RAND_3271;
  reg [31:0] _RAND_3272;
  reg [31:0] _RAND_3273;
  reg [31:0] _RAND_3274;
  reg [31:0] _RAND_3275;
  reg [31:0] _RAND_3276;
  reg [31:0] _RAND_3277;
  reg [31:0] _RAND_3278;
  reg [31:0] _RAND_3279;
  reg [31:0] _RAND_3280;
  reg [31:0] _RAND_3281;
  reg [31:0] _RAND_3282;
  reg [31:0] _RAND_3283;
  reg [31:0] _RAND_3284;
  reg [31:0] _RAND_3285;
  reg [31:0] _RAND_3286;
  reg [31:0] _RAND_3287;
  reg [31:0] _RAND_3288;
  reg [31:0] _RAND_3289;
  reg [31:0] _RAND_3290;
  reg [31:0] _RAND_3291;
  reg [31:0] _RAND_3292;
  reg [31:0] _RAND_3293;
  reg [31:0] _RAND_3294;
  reg [31:0] _RAND_3295;
  reg [31:0] _RAND_3296;
  reg [31:0] _RAND_3297;
  reg [31:0] _RAND_3298;
  reg [31:0] _RAND_3299;
  reg [31:0] _RAND_3300;
  reg [31:0] _RAND_3301;
  reg [31:0] _RAND_3302;
  reg [31:0] _RAND_3303;
  reg [31:0] _RAND_3304;
  reg [31:0] _RAND_3305;
  reg [31:0] _RAND_3306;
  reg [31:0] _RAND_3307;
  reg [31:0] _RAND_3308;
  reg [31:0] _RAND_3309;
  reg [31:0] _RAND_3310;
  reg [31:0] _RAND_3311;
  reg [31:0] _RAND_3312;
  reg [31:0] _RAND_3313;
  reg [31:0] _RAND_3314;
  reg [31:0] _RAND_3315;
  reg [31:0] _RAND_3316;
  reg [31:0] _RAND_3317;
  reg [31:0] _RAND_3318;
  reg [31:0] _RAND_3319;
  reg [31:0] _RAND_3320;
  reg [31:0] _RAND_3321;
  reg [31:0] _RAND_3322;
  reg [31:0] _RAND_3323;
  reg [31:0] _RAND_3324;
  reg [31:0] _RAND_3325;
  reg [31:0] _RAND_3326;
  reg [31:0] _RAND_3327;
  reg [31:0] _RAND_3328;
  reg [31:0] _RAND_3329;
  reg [31:0] _RAND_3330;
  reg [31:0] _RAND_3331;
  reg [31:0] _RAND_3332;
  reg [31:0] _RAND_3333;
  reg [31:0] _RAND_3334;
  reg [31:0] _RAND_3335;
  reg [31:0] _RAND_3336;
  reg [31:0] _RAND_3337;
  reg [31:0] _RAND_3338;
  reg [31:0] _RAND_3339;
  reg [31:0] _RAND_3340;
  reg [31:0] _RAND_3341;
  reg [31:0] _RAND_3342;
  reg [31:0] _RAND_3343;
  reg [31:0] _RAND_3344;
  reg [31:0] _RAND_3345;
  reg [31:0] _RAND_3346;
  reg [31:0] _RAND_3347;
  reg [31:0] _RAND_3348;
  reg [31:0] _RAND_3349;
  reg [31:0] _RAND_3350;
  reg [31:0] _RAND_3351;
  reg [31:0] _RAND_3352;
  reg [31:0] _RAND_3353;
  reg [31:0] _RAND_3354;
  reg [31:0] _RAND_3355;
  reg [31:0] _RAND_3356;
  reg [31:0] _RAND_3357;
  reg [31:0] _RAND_3358;
  reg [31:0] _RAND_3359;
  reg [31:0] _RAND_3360;
  reg [31:0] _RAND_3361;
  reg [31:0] _RAND_3362;
  reg [31:0] _RAND_3363;
  reg [31:0] _RAND_3364;
  reg [31:0] _RAND_3365;
  reg [31:0] _RAND_3366;
  reg [31:0] _RAND_3367;
  reg [31:0] _RAND_3368;
  reg [31:0] _RAND_3369;
  reg [31:0] _RAND_3370;
  reg [31:0] _RAND_3371;
  reg [31:0] _RAND_3372;
  reg [31:0] _RAND_3373;
  reg [31:0] _RAND_3374;
  reg [31:0] _RAND_3375;
  reg [31:0] _RAND_3376;
  reg [31:0] _RAND_3377;
  reg [31:0] _RAND_3378;
  reg [31:0] _RAND_3379;
  reg [31:0] _RAND_3380;
  reg [31:0] _RAND_3381;
  reg [31:0] _RAND_3382;
  reg [31:0] _RAND_3383;
  reg [31:0] _RAND_3384;
  reg [31:0] _RAND_3385;
  reg [31:0] _RAND_3386;
  reg [31:0] _RAND_3387;
  reg [31:0] _RAND_3388;
  reg [31:0] _RAND_3389;
  reg [31:0] _RAND_3390;
  reg [31:0] _RAND_3391;
  reg [31:0] _RAND_3392;
  reg [31:0] _RAND_3393;
  reg [31:0] _RAND_3394;
  reg [31:0] _RAND_3395;
  reg [31:0] _RAND_3396;
  reg [31:0] _RAND_3397;
  reg [31:0] _RAND_3398;
  reg [31:0] _RAND_3399;
  reg [31:0] _RAND_3400;
  reg [31:0] _RAND_3401;
  reg [31:0] _RAND_3402;
  reg [31:0] _RAND_3403;
  reg [31:0] _RAND_3404;
  reg [31:0] _RAND_3405;
  reg [31:0] _RAND_3406;
  reg [31:0] _RAND_3407;
  reg [31:0] _RAND_3408;
  reg [31:0] _RAND_3409;
  reg [31:0] _RAND_3410;
  reg [31:0] _RAND_3411;
  reg [31:0] _RAND_3412;
  reg [31:0] _RAND_3413;
  reg [31:0] _RAND_3414;
  reg [31:0] _RAND_3415;
  reg [31:0] _RAND_3416;
  reg [31:0] _RAND_3417;
  reg [31:0] _RAND_3418;
  reg [31:0] _RAND_3419;
  reg [31:0] _RAND_3420;
  reg [31:0] _RAND_3421;
  reg [31:0] _RAND_3422;
  reg [31:0] _RAND_3423;
  reg [31:0] _RAND_3424;
  reg [31:0] _RAND_3425;
  reg [31:0] _RAND_3426;
  reg [31:0] _RAND_3427;
  reg [31:0] _RAND_3428;
  reg [31:0] _RAND_3429;
  reg [31:0] _RAND_3430;
  reg [31:0] _RAND_3431;
  reg [31:0] _RAND_3432;
  reg [31:0] _RAND_3433;
  reg [31:0] _RAND_3434;
  reg [31:0] _RAND_3435;
  reg [31:0] _RAND_3436;
  reg [31:0] _RAND_3437;
  reg [31:0] _RAND_3438;
  reg [31:0] _RAND_3439;
  reg [31:0] _RAND_3440;
  reg [31:0] _RAND_3441;
  reg [31:0] _RAND_3442;
  reg [31:0] _RAND_3443;
  reg [31:0] _RAND_3444;
  reg [31:0] _RAND_3445;
  reg [31:0] _RAND_3446;
  reg [31:0] _RAND_3447;
  reg [31:0] _RAND_3448;
  reg [31:0] _RAND_3449;
  reg [31:0] _RAND_3450;
  reg [31:0] _RAND_3451;
  reg [31:0] _RAND_3452;
  reg [31:0] _RAND_3453;
  reg [31:0] _RAND_3454;
  reg [31:0] _RAND_3455;
  reg [31:0] _RAND_3456;
  reg [31:0] _RAND_3457;
  reg [31:0] _RAND_3458;
  reg [31:0] _RAND_3459;
  reg [31:0] _RAND_3460;
  reg [31:0] _RAND_3461;
  reg [31:0] _RAND_3462;
  reg [31:0] _RAND_3463;
  reg [31:0] _RAND_3464;
  reg [31:0] _RAND_3465;
  reg [31:0] _RAND_3466;
  reg [31:0] _RAND_3467;
  reg [31:0] _RAND_3468;
  reg [31:0] _RAND_3469;
  reg [31:0] _RAND_3470;
  reg [31:0] _RAND_3471;
  reg [31:0] _RAND_3472;
  reg [31:0] _RAND_3473;
  reg [31:0] _RAND_3474;
  reg [31:0] _RAND_3475;
  reg [31:0] _RAND_3476;
  reg [31:0] _RAND_3477;
  reg [31:0] _RAND_3478;
  reg [31:0] _RAND_3479;
  reg [31:0] _RAND_3480;
  reg [31:0] _RAND_3481;
  reg [31:0] _RAND_3482;
  reg [31:0] _RAND_3483;
  reg [31:0] _RAND_3484;
  reg [31:0] _RAND_3485;
  reg [31:0] _RAND_3486;
  reg [31:0] _RAND_3487;
  reg [31:0] _RAND_3488;
  reg [31:0] _RAND_3489;
  reg [31:0] _RAND_3490;
  reg [31:0] _RAND_3491;
  reg [31:0] _RAND_3492;
  reg [31:0] _RAND_3493;
  reg [31:0] _RAND_3494;
  reg [31:0] _RAND_3495;
  reg [31:0] _RAND_3496;
  reg [31:0] _RAND_3497;
  reg [31:0] _RAND_3498;
  reg [31:0] _RAND_3499;
  reg [31:0] _RAND_3500;
  reg [31:0] _RAND_3501;
  reg [31:0] _RAND_3502;
  reg [31:0] _RAND_3503;
  reg [31:0] _RAND_3504;
  reg [31:0] _RAND_3505;
  reg [31:0] _RAND_3506;
  reg [31:0] _RAND_3507;
  reg [31:0] _RAND_3508;
  reg [31:0] _RAND_3509;
  reg [31:0] _RAND_3510;
  reg [31:0] _RAND_3511;
  reg [31:0] _RAND_3512;
  reg [31:0] _RAND_3513;
  reg [31:0] _RAND_3514;
  reg [31:0] _RAND_3515;
  reg [31:0] _RAND_3516;
  reg [31:0] _RAND_3517;
  reg [31:0] _RAND_3518;
  reg [31:0] _RAND_3519;
  reg [31:0] _RAND_3520;
  reg [31:0] _RAND_3521;
  reg [31:0] _RAND_3522;
  reg [31:0] _RAND_3523;
  reg [31:0] _RAND_3524;
  reg [31:0] _RAND_3525;
  reg [31:0] _RAND_3526;
  reg [31:0] _RAND_3527;
  reg [31:0] _RAND_3528;
  reg [31:0] _RAND_3529;
  reg [31:0] _RAND_3530;
  reg [31:0] _RAND_3531;
  reg [31:0] _RAND_3532;
  reg [31:0] _RAND_3533;
  reg [31:0] _RAND_3534;
  reg [31:0] _RAND_3535;
  reg [31:0] _RAND_3536;
  reg [31:0] _RAND_3537;
  reg [31:0] _RAND_3538;
  reg [31:0] _RAND_3539;
  reg [31:0] _RAND_3540;
  reg [31:0] _RAND_3541;
  reg [31:0] _RAND_3542;
  reg [31:0] _RAND_3543;
  reg [31:0] _RAND_3544;
  reg [31:0] _RAND_3545;
  reg [31:0] _RAND_3546;
  reg [31:0] _RAND_3547;
  reg [31:0] _RAND_3548;
  reg [31:0] _RAND_3549;
  reg [31:0] _RAND_3550;
  reg [31:0] _RAND_3551;
  reg [31:0] _RAND_3552;
  reg [31:0] _RAND_3553;
  reg [31:0] _RAND_3554;
  reg [31:0] _RAND_3555;
  reg [31:0] _RAND_3556;
  reg [31:0] _RAND_3557;
  reg [31:0] _RAND_3558;
  reg [31:0] _RAND_3559;
  reg [31:0] _RAND_3560;
  reg [31:0] _RAND_3561;
  reg [31:0] _RAND_3562;
  reg [31:0] _RAND_3563;
  reg [31:0] _RAND_3564;
  reg [31:0] _RAND_3565;
  reg [31:0] _RAND_3566;
  reg [31:0] _RAND_3567;
  reg [31:0] _RAND_3568;
  reg [31:0] _RAND_3569;
  reg [31:0] _RAND_3570;
  reg [31:0] _RAND_3571;
  reg [31:0] _RAND_3572;
  reg [31:0] _RAND_3573;
  reg [31:0] _RAND_3574;
  reg [31:0] _RAND_3575;
  reg [31:0] _RAND_3576;
  reg [31:0] _RAND_3577;
  reg [31:0] _RAND_3578;
  reg [31:0] _RAND_3579;
  reg [31:0] _RAND_3580;
  reg [31:0] _RAND_3581;
  reg [31:0] _RAND_3582;
  reg [31:0] _RAND_3583;
  reg [31:0] _RAND_3584;
  reg [31:0] _RAND_3585;
  reg [31:0] _RAND_3586;
  reg [31:0] _RAND_3587;
  reg [31:0] _RAND_3588;
  reg [31:0] _RAND_3589;
  reg [31:0] _RAND_3590;
  reg [31:0] _RAND_3591;
  reg [31:0] _RAND_3592;
  reg [31:0] _RAND_3593;
  reg [31:0] _RAND_3594;
  reg [31:0] _RAND_3595;
  reg [31:0] _RAND_3596;
  reg [31:0] _RAND_3597;
  reg [31:0] _RAND_3598;
  reg [31:0] _RAND_3599;
  reg [31:0] _RAND_3600;
  reg [31:0] _RAND_3601;
  reg [31:0] _RAND_3602;
  reg [31:0] _RAND_3603;
  reg [31:0] _RAND_3604;
  reg [31:0] _RAND_3605;
  reg [31:0] _RAND_3606;
  reg [31:0] _RAND_3607;
  reg [31:0] _RAND_3608;
  reg [31:0] _RAND_3609;
  reg [31:0] _RAND_3610;
  reg [31:0] _RAND_3611;
  reg [31:0] _RAND_3612;
  reg [31:0] _RAND_3613;
  reg [31:0] _RAND_3614;
  reg [31:0] _RAND_3615;
  reg [31:0] _RAND_3616;
  reg [31:0] _RAND_3617;
  reg [31:0] _RAND_3618;
  reg [31:0] _RAND_3619;
  reg [31:0] _RAND_3620;
  reg [31:0] _RAND_3621;
  reg [31:0] _RAND_3622;
  reg [31:0] _RAND_3623;
  reg [31:0] _RAND_3624;
  reg [31:0] _RAND_3625;
  reg [31:0] _RAND_3626;
  reg [31:0] _RAND_3627;
  reg [31:0] _RAND_3628;
  reg [31:0] _RAND_3629;
  reg [31:0] _RAND_3630;
  reg [31:0] _RAND_3631;
  reg [31:0] _RAND_3632;
  reg [31:0] _RAND_3633;
  reg [31:0] _RAND_3634;
  reg [31:0] _RAND_3635;
  reg [31:0] _RAND_3636;
  reg [31:0] _RAND_3637;
  reg [31:0] _RAND_3638;
  reg [31:0] _RAND_3639;
  reg [31:0] _RAND_3640;
  reg [31:0] _RAND_3641;
  reg [31:0] _RAND_3642;
  reg [31:0] _RAND_3643;
  reg [31:0] _RAND_3644;
  reg [31:0] _RAND_3645;
  reg [31:0] _RAND_3646;
  reg [31:0] _RAND_3647;
  reg [31:0] _RAND_3648;
  reg [31:0] _RAND_3649;
  reg [31:0] _RAND_3650;
  reg [31:0] _RAND_3651;
  reg [31:0] _RAND_3652;
  reg [31:0] _RAND_3653;
  reg [31:0] _RAND_3654;
  reg [31:0] _RAND_3655;
  reg [31:0] _RAND_3656;
  reg [31:0] _RAND_3657;
  reg [31:0] _RAND_3658;
  reg [31:0] _RAND_3659;
  reg [31:0] _RAND_3660;
  reg [31:0] _RAND_3661;
  reg [31:0] _RAND_3662;
  reg [31:0] _RAND_3663;
  reg [31:0] _RAND_3664;
  reg [31:0] _RAND_3665;
  reg [31:0] _RAND_3666;
  reg [31:0] _RAND_3667;
  reg [31:0] _RAND_3668;
  reg [31:0] _RAND_3669;
  reg [31:0] _RAND_3670;
  reg [31:0] _RAND_3671;
  reg [31:0] _RAND_3672;
  reg [31:0] _RAND_3673;
  reg [31:0] _RAND_3674;
  reg [31:0] _RAND_3675;
  reg [31:0] _RAND_3676;
  reg [31:0] _RAND_3677;
  reg [31:0] _RAND_3678;
  reg [31:0] _RAND_3679;
  reg [31:0] _RAND_3680;
  reg [31:0] _RAND_3681;
  reg [31:0] _RAND_3682;
  reg [31:0] _RAND_3683;
  reg [31:0] _RAND_3684;
  reg [31:0] _RAND_3685;
  reg [31:0] _RAND_3686;
  reg [31:0] _RAND_3687;
  reg [31:0] _RAND_3688;
  reg [31:0] _RAND_3689;
  reg [31:0] _RAND_3690;
  reg [31:0] _RAND_3691;
  reg [31:0] _RAND_3692;
  reg [31:0] _RAND_3693;
  reg [31:0] _RAND_3694;
  reg [31:0] _RAND_3695;
  reg [31:0] _RAND_3696;
  reg [31:0] _RAND_3697;
  reg [31:0] _RAND_3698;
  reg [31:0] _RAND_3699;
  reg [31:0] _RAND_3700;
  reg [31:0] _RAND_3701;
  reg [31:0] _RAND_3702;
  reg [31:0] _RAND_3703;
  reg [31:0] _RAND_3704;
  reg [31:0] _RAND_3705;
  reg [31:0] _RAND_3706;
  reg [31:0] _RAND_3707;
  reg [31:0] _RAND_3708;
  reg [31:0] _RAND_3709;
  reg [31:0] _RAND_3710;
  reg [31:0] _RAND_3711;
  reg [31:0] _RAND_3712;
  reg [31:0] _RAND_3713;
  reg [31:0] _RAND_3714;
  reg [31:0] _RAND_3715;
  reg [31:0] _RAND_3716;
  reg [31:0] _RAND_3717;
  reg [31:0] _RAND_3718;
  reg [31:0] _RAND_3719;
  reg [31:0] _RAND_3720;
  reg [31:0] _RAND_3721;
  reg [31:0] _RAND_3722;
  reg [31:0] _RAND_3723;
  reg [31:0] _RAND_3724;
  reg [31:0] _RAND_3725;
  reg [31:0] _RAND_3726;
  reg [31:0] _RAND_3727;
  reg [31:0] _RAND_3728;
  reg [31:0] _RAND_3729;
  reg [31:0] _RAND_3730;
  reg [31:0] _RAND_3731;
  reg [31:0] _RAND_3732;
  reg [31:0] _RAND_3733;
  reg [31:0] _RAND_3734;
  reg [31:0] _RAND_3735;
  reg [31:0] _RAND_3736;
  reg [31:0] _RAND_3737;
  reg [31:0] _RAND_3738;
  reg [31:0] _RAND_3739;
  reg [31:0] _RAND_3740;
  reg [31:0] _RAND_3741;
  reg [31:0] _RAND_3742;
  reg [31:0] _RAND_3743;
  reg [31:0] _RAND_3744;
  reg [31:0] _RAND_3745;
  reg [31:0] _RAND_3746;
  reg [31:0] _RAND_3747;
  reg [31:0] _RAND_3748;
  reg [31:0] _RAND_3749;
  reg [31:0] _RAND_3750;
  reg [31:0] _RAND_3751;
  reg [31:0] _RAND_3752;
  reg [31:0] _RAND_3753;
  reg [31:0] _RAND_3754;
  reg [31:0] _RAND_3755;
  reg [31:0] _RAND_3756;
  reg [31:0] _RAND_3757;
  reg [31:0] _RAND_3758;
  reg [31:0] _RAND_3759;
  reg [31:0] _RAND_3760;
  reg [31:0] _RAND_3761;
  reg [31:0] _RAND_3762;
  reg [31:0] _RAND_3763;
  reg [31:0] _RAND_3764;
  reg [31:0] _RAND_3765;
  reg [31:0] _RAND_3766;
  reg [31:0] _RAND_3767;
  reg [31:0] _RAND_3768;
  reg [31:0] _RAND_3769;
  reg [31:0] _RAND_3770;
  reg [31:0] _RAND_3771;
  reg [31:0] _RAND_3772;
  reg [31:0] _RAND_3773;
  reg [31:0] _RAND_3774;
  reg [31:0] _RAND_3775;
  reg [31:0] _RAND_3776;
  reg [31:0] _RAND_3777;
  reg [31:0] _RAND_3778;
  reg [31:0] _RAND_3779;
  reg [31:0] _RAND_3780;
  reg [31:0] _RAND_3781;
  reg [31:0] _RAND_3782;
  reg [31:0] _RAND_3783;
  reg [31:0] _RAND_3784;
  reg [31:0] _RAND_3785;
  reg [31:0] _RAND_3786;
  reg [31:0] _RAND_3787;
  reg [31:0] _RAND_3788;
  reg [31:0] _RAND_3789;
  reg [31:0] _RAND_3790;
  reg [31:0] _RAND_3791;
  reg [31:0] _RAND_3792;
  reg [31:0] _RAND_3793;
  reg [31:0] _RAND_3794;
  reg [31:0] _RAND_3795;
  reg [31:0] _RAND_3796;
  reg [31:0] _RAND_3797;
  reg [31:0] _RAND_3798;
  reg [31:0] _RAND_3799;
  reg [31:0] _RAND_3800;
  reg [31:0] _RAND_3801;
  reg [31:0] _RAND_3802;
  reg [31:0] _RAND_3803;
  reg [31:0] _RAND_3804;
  reg [31:0] _RAND_3805;
  reg [31:0] _RAND_3806;
  reg [31:0] _RAND_3807;
  reg [31:0] _RAND_3808;
  reg [31:0] _RAND_3809;
  reg [31:0] _RAND_3810;
  reg [31:0] _RAND_3811;
  reg [31:0] _RAND_3812;
  reg [31:0] _RAND_3813;
  reg [31:0] _RAND_3814;
  reg [31:0] _RAND_3815;
  reg [31:0] _RAND_3816;
  reg [31:0] _RAND_3817;
  reg [31:0] _RAND_3818;
  reg [31:0] _RAND_3819;
  reg [31:0] _RAND_3820;
  reg [31:0] _RAND_3821;
  reg [31:0] _RAND_3822;
  reg [31:0] _RAND_3823;
  reg [31:0] _RAND_3824;
  reg [31:0] _RAND_3825;
  reg [31:0] _RAND_3826;
  reg [31:0] _RAND_3827;
  reg [31:0] _RAND_3828;
  reg [31:0] _RAND_3829;
  reg [31:0] _RAND_3830;
  reg [31:0] _RAND_3831;
  reg [31:0] _RAND_3832;
  reg [31:0] _RAND_3833;
  reg [31:0] _RAND_3834;
  reg [31:0] _RAND_3835;
  reg [31:0] _RAND_3836;
  reg [31:0] _RAND_3837;
  reg [31:0] _RAND_3838;
  reg [31:0] _RAND_3839;
  reg [31:0] _RAND_3840;
  reg [31:0] _RAND_3841;
  reg [31:0] _RAND_3842;
  reg [31:0] _RAND_3843;
  reg [31:0] _RAND_3844;
  reg [31:0] _RAND_3845;
  reg [31:0] _RAND_3846;
  reg [31:0] _RAND_3847;
  reg [31:0] _RAND_3848;
  reg [31:0] _RAND_3849;
  reg [31:0] _RAND_3850;
  reg [31:0] _RAND_3851;
  reg [31:0] _RAND_3852;
  reg [31:0] _RAND_3853;
  reg [31:0] _RAND_3854;
  reg [31:0] _RAND_3855;
  reg [31:0] _RAND_3856;
  reg [31:0] _RAND_3857;
  reg [31:0] _RAND_3858;
  reg [31:0] _RAND_3859;
  reg [31:0] _RAND_3860;
  reg [31:0] _RAND_3861;
  reg [31:0] _RAND_3862;
  reg [31:0] _RAND_3863;
  reg [31:0] _RAND_3864;
  reg [31:0] _RAND_3865;
  reg [31:0] _RAND_3866;
  reg [31:0] _RAND_3867;
  reg [31:0] _RAND_3868;
  reg [31:0] _RAND_3869;
  reg [31:0] _RAND_3870;
  reg [31:0] _RAND_3871;
  reg [31:0] _RAND_3872;
  reg [31:0] _RAND_3873;
  reg [31:0] _RAND_3874;
  reg [31:0] _RAND_3875;
  reg [31:0] _RAND_3876;
  reg [31:0] _RAND_3877;
  reg [31:0] _RAND_3878;
  reg [31:0] _RAND_3879;
  reg [31:0] _RAND_3880;
  reg [31:0] _RAND_3881;
  reg [31:0] _RAND_3882;
  reg [31:0] _RAND_3883;
  reg [31:0] _RAND_3884;
  reg [31:0] _RAND_3885;
  reg [31:0] _RAND_3886;
  reg [31:0] _RAND_3887;
  reg [31:0] _RAND_3888;
  reg [31:0] _RAND_3889;
  reg [31:0] _RAND_3890;
  reg [31:0] _RAND_3891;
  reg [31:0] _RAND_3892;
  reg [31:0] _RAND_3893;
  reg [31:0] _RAND_3894;
  reg [31:0] _RAND_3895;
  reg [31:0] _RAND_3896;
  reg [31:0] _RAND_3897;
  reg [31:0] _RAND_3898;
  reg [31:0] _RAND_3899;
  reg [31:0] _RAND_3900;
  reg [31:0] _RAND_3901;
  reg [31:0] _RAND_3902;
  reg [31:0] _RAND_3903;
  reg [31:0] _RAND_3904;
  reg [31:0] _RAND_3905;
  reg [31:0] _RAND_3906;
  reg [31:0] _RAND_3907;
  reg [31:0] _RAND_3908;
  reg [31:0] _RAND_3909;
  reg [31:0] _RAND_3910;
  reg [31:0] _RAND_3911;
  reg [31:0] _RAND_3912;
  reg [31:0] _RAND_3913;
  reg [31:0] _RAND_3914;
  reg [31:0] _RAND_3915;
  reg [31:0] _RAND_3916;
  reg [31:0] _RAND_3917;
  reg [31:0] _RAND_3918;
  reg [31:0] _RAND_3919;
  reg [31:0] _RAND_3920;
  reg [31:0] _RAND_3921;
  reg [31:0] _RAND_3922;
  reg [31:0] _RAND_3923;
  reg [31:0] _RAND_3924;
  reg [31:0] _RAND_3925;
  reg [31:0] _RAND_3926;
  reg [31:0] _RAND_3927;
  reg [31:0] _RAND_3928;
  reg [31:0] _RAND_3929;
  reg [31:0] _RAND_3930;
  reg [31:0] _RAND_3931;
  reg [31:0] _RAND_3932;
  reg [31:0] _RAND_3933;
  reg [31:0] _RAND_3934;
  reg [31:0] _RAND_3935;
  reg [31:0] _RAND_3936;
  reg [31:0] _RAND_3937;
  reg [31:0] _RAND_3938;
  reg [31:0] _RAND_3939;
  reg [31:0] _RAND_3940;
  reg [31:0] _RAND_3941;
  reg [31:0] _RAND_3942;
  reg [31:0] _RAND_3943;
  reg [31:0] _RAND_3944;
  reg [31:0] _RAND_3945;
  reg [31:0] _RAND_3946;
  reg [31:0] _RAND_3947;
  reg [31:0] _RAND_3948;
  reg [31:0] _RAND_3949;
  reg [31:0] _RAND_3950;
  reg [31:0] _RAND_3951;
  reg [31:0] _RAND_3952;
  reg [31:0] _RAND_3953;
  reg [31:0] _RAND_3954;
  reg [31:0] _RAND_3955;
  reg [31:0] _RAND_3956;
  reg [31:0] _RAND_3957;
  reg [31:0] _RAND_3958;
  reg [31:0] _RAND_3959;
  reg [31:0] _RAND_3960;
  reg [31:0] _RAND_3961;
  reg [31:0] _RAND_3962;
  reg [31:0] _RAND_3963;
  reg [31:0] _RAND_3964;
  reg [31:0] _RAND_3965;
  reg [31:0] _RAND_3966;
  reg [31:0] _RAND_3967;
  reg [31:0] _RAND_3968;
  reg [31:0] _RAND_3969;
  reg [31:0] _RAND_3970;
  reg [31:0] _RAND_3971;
  reg [31:0] _RAND_3972;
  reg [31:0] _RAND_3973;
  reg [31:0] _RAND_3974;
  reg [31:0] _RAND_3975;
  reg [31:0] _RAND_3976;
  reg [31:0] _RAND_3977;
  reg [31:0] _RAND_3978;
  reg [31:0] _RAND_3979;
  reg [31:0] _RAND_3980;
  reg [31:0] _RAND_3981;
  reg [31:0] _RAND_3982;
  reg [31:0] _RAND_3983;
  reg [31:0] _RAND_3984;
  reg [31:0] _RAND_3985;
  reg [31:0] _RAND_3986;
  reg [31:0] _RAND_3987;
  reg [31:0] _RAND_3988;
  reg [31:0] _RAND_3989;
  reg [31:0] _RAND_3990;
  reg [31:0] _RAND_3991;
  reg [31:0] _RAND_3992;
  reg [31:0] _RAND_3993;
  reg [31:0] _RAND_3994;
  reg [31:0] _RAND_3995;
  reg [31:0] _RAND_3996;
  reg [31:0] _RAND_3997;
  reg [31:0] _RAND_3998;
  reg [31:0] _RAND_3999;
  reg [31:0] _RAND_4000;
  reg [31:0] _RAND_4001;
  reg [31:0] _RAND_4002;
  reg [31:0] _RAND_4003;
  reg [31:0] _RAND_4004;
  reg [31:0] _RAND_4005;
  reg [31:0] _RAND_4006;
  reg [31:0] _RAND_4007;
  reg [31:0] _RAND_4008;
  reg [31:0] _RAND_4009;
  reg [31:0] _RAND_4010;
  reg [31:0] _RAND_4011;
  reg [31:0] _RAND_4012;
  reg [31:0] _RAND_4013;
  reg [31:0] _RAND_4014;
  reg [31:0] _RAND_4015;
  reg [31:0] _RAND_4016;
  reg [31:0] _RAND_4017;
  reg [31:0] _RAND_4018;
  reg [31:0] _RAND_4019;
  reg [31:0] _RAND_4020;
  reg [31:0] _RAND_4021;
  reg [31:0] _RAND_4022;
  reg [31:0] _RAND_4023;
  reg [31:0] _RAND_4024;
  reg [31:0] _RAND_4025;
  reg [31:0] _RAND_4026;
  reg [31:0] _RAND_4027;
  reg [31:0] _RAND_4028;
  reg [31:0] _RAND_4029;
  reg [31:0] _RAND_4030;
  reg [31:0] _RAND_4031;
  reg [31:0] _RAND_4032;
  reg [31:0] _RAND_4033;
  reg [31:0] _RAND_4034;
  reg [31:0] _RAND_4035;
  reg [31:0] _RAND_4036;
  reg [31:0] _RAND_4037;
  reg [31:0] _RAND_4038;
  reg [31:0] _RAND_4039;
  reg [31:0] _RAND_4040;
  reg [31:0] _RAND_4041;
  reg [31:0] _RAND_4042;
  reg [31:0] _RAND_4043;
  reg [31:0] _RAND_4044;
  reg [31:0] _RAND_4045;
  reg [31:0] _RAND_4046;
  reg [31:0] _RAND_4047;
  reg [31:0] _RAND_4048;
  reg [31:0] _RAND_4049;
  reg [31:0] _RAND_4050;
  reg [31:0] _RAND_4051;
  reg [31:0] _RAND_4052;
  reg [31:0] _RAND_4053;
  reg [31:0] _RAND_4054;
  reg [31:0] _RAND_4055;
  reg [31:0] _RAND_4056;
  reg [31:0] _RAND_4057;
  reg [31:0] _RAND_4058;
  reg [31:0] _RAND_4059;
  reg [31:0] _RAND_4060;
  reg [31:0] _RAND_4061;
  reg [31:0] _RAND_4062;
  reg [31:0] _RAND_4063;
  reg [31:0] _RAND_4064;
  reg [31:0] _RAND_4065;
  reg [31:0] _RAND_4066;
  reg [31:0] _RAND_4067;
  reg [31:0] _RAND_4068;
  reg [31:0] _RAND_4069;
  reg [31:0] _RAND_4070;
  reg [31:0] _RAND_4071;
  reg [31:0] _RAND_4072;
  reg [31:0] _RAND_4073;
  reg [31:0] _RAND_4074;
  reg [31:0] _RAND_4075;
  reg [31:0] _RAND_4076;
  reg [31:0] _RAND_4077;
  reg [31:0] _RAND_4078;
  reg [31:0] _RAND_4079;
  reg [31:0] _RAND_4080;
  reg [31:0] _RAND_4081;
  reg [31:0] _RAND_4082;
  reg [31:0] _RAND_4083;
  reg [31:0] _RAND_4084;
  reg [31:0] _RAND_4085;
  reg [31:0] _RAND_4086;
  reg [31:0] _RAND_4087;
  reg [31:0] _RAND_4088;
  reg [31:0] _RAND_4089;
  reg [31:0] _RAND_4090;
  reg [31:0] _RAND_4091;
  reg [31:0] _RAND_4092;
  reg [31:0] _RAND_4093;
  reg [31:0] _RAND_4094;
  reg [31:0] _RAND_4095;
  reg [31:0] _RAND_4096;
  reg [31:0] _RAND_4097;
  reg [31:0] _RAND_4098;
  reg [31:0] _RAND_4099;
  reg [31:0] _RAND_4100;
  reg [31:0] _RAND_4101;
  reg [31:0] _RAND_4102;
  reg [31:0] _RAND_4103;
  reg [31:0] _RAND_4104;
  reg [31:0] _RAND_4105;
  reg [31:0] _RAND_4106;
  reg [31:0] _RAND_4107;
  reg [31:0] _RAND_4108;
  reg [31:0] _RAND_4109;
  reg [31:0] _RAND_4110;
  reg [31:0] _RAND_4111;
  reg [31:0] _RAND_4112;
  reg [31:0] _RAND_4113;
  reg [31:0] _RAND_4114;
  reg [31:0] _RAND_4115;
  reg [31:0] _RAND_4116;
  reg [31:0] _RAND_4117;
  reg [31:0] _RAND_4118;
  reg [31:0] _RAND_4119;
  reg [31:0] _RAND_4120;
  reg [31:0] _RAND_4121;
  reg [31:0] _RAND_4122;
  reg [31:0] _RAND_4123;
  reg [31:0] _RAND_4124;
  reg [31:0] _RAND_4125;
  reg [31:0] _RAND_4126;
  reg [31:0] _RAND_4127;
  reg [31:0] _RAND_4128;
  reg [31:0] _RAND_4129;
  reg [31:0] _RAND_4130;
  reg [31:0] _RAND_4131;
  reg [31:0] _RAND_4132;
  reg [31:0] _RAND_4133;
  reg [31:0] _RAND_4134;
  reg [31:0] _RAND_4135;
  reg [31:0] _RAND_4136;
  reg [31:0] _RAND_4137;
  reg [31:0] _RAND_4138;
  reg [31:0] _RAND_4139;
  reg [31:0] _RAND_4140;
  reg [31:0] _RAND_4141;
  reg [31:0] _RAND_4142;
  reg [31:0] _RAND_4143;
  reg [31:0] _RAND_4144;
  reg [31:0] _RAND_4145;
  reg [31:0] _RAND_4146;
  reg [31:0] _RAND_4147;
  reg [31:0] _RAND_4148;
  reg [31:0] _RAND_4149;
  reg [31:0] _RAND_4150;
  reg [31:0] _RAND_4151;
  reg [31:0] _RAND_4152;
  reg [31:0] _RAND_4153;
  reg [31:0] _RAND_4154;
  reg [31:0] _RAND_4155;
  reg [31:0] _RAND_4156;
  reg [31:0] _RAND_4157;
  reg [31:0] _RAND_4158;
  reg [31:0] _RAND_4159;
  reg [31:0] _RAND_4160;
  reg [31:0] _RAND_4161;
  reg [31:0] _RAND_4162;
  reg [31:0] _RAND_4163;
  reg [31:0] _RAND_4164;
  reg [31:0] _RAND_4165;
  reg [31:0] _RAND_4166;
  reg [31:0] _RAND_4167;
  reg [31:0] _RAND_4168;
  reg [31:0] _RAND_4169;
  reg [31:0] _RAND_4170;
  reg [31:0] _RAND_4171;
  reg [31:0] _RAND_4172;
  reg [31:0] _RAND_4173;
  reg [31:0] _RAND_4174;
  reg [31:0] _RAND_4175;
  reg [31:0] _RAND_4176;
  reg [31:0] _RAND_4177;
  reg [31:0] _RAND_4178;
  reg [31:0] _RAND_4179;
  reg [31:0] _RAND_4180;
  reg [31:0] _RAND_4181;
  reg [31:0] _RAND_4182;
  reg [31:0] _RAND_4183;
  reg [31:0] _RAND_4184;
  reg [31:0] _RAND_4185;
  reg [31:0] _RAND_4186;
  reg [31:0] _RAND_4187;
  reg [31:0] _RAND_4188;
  reg [31:0] _RAND_4189;
  reg [31:0] _RAND_4190;
  reg [31:0] _RAND_4191;
  reg [31:0] _RAND_4192;
  reg [31:0] _RAND_4193;
  reg [31:0] _RAND_4194;
  reg [31:0] _RAND_4195;
  reg [31:0] _RAND_4196;
  reg [31:0] _RAND_4197;
  reg [31:0] _RAND_4198;
  reg [31:0] _RAND_4199;
  reg [31:0] _RAND_4200;
  reg [31:0] _RAND_4201;
  reg [31:0] _RAND_4202;
  reg [31:0] _RAND_4203;
  reg [31:0] _RAND_4204;
  reg [31:0] _RAND_4205;
  reg [31:0] _RAND_4206;
  reg [31:0] _RAND_4207;
  reg [31:0] _RAND_4208;
  reg [31:0] _RAND_4209;
  reg [31:0] _RAND_4210;
  reg [31:0] _RAND_4211;
  reg [31:0] _RAND_4212;
  reg [31:0] _RAND_4213;
  reg [31:0] _RAND_4214;
  reg [31:0] _RAND_4215;
  reg [31:0] _RAND_4216;
  reg [31:0] _RAND_4217;
  reg [31:0] _RAND_4218;
  reg [31:0] _RAND_4219;
  reg [31:0] _RAND_4220;
  reg [31:0] _RAND_4221;
  reg [31:0] _RAND_4222;
  reg [31:0] _RAND_4223;
  reg [31:0] _RAND_4224;
  reg [31:0] _RAND_4225;
  reg [31:0] _RAND_4226;
  reg [31:0] _RAND_4227;
  reg [31:0] _RAND_4228;
  reg [31:0] _RAND_4229;
  reg [31:0] _RAND_4230;
  reg [31:0] _RAND_4231;
  reg [31:0] _RAND_4232;
  reg [31:0] _RAND_4233;
  reg [31:0] _RAND_4234;
  reg [31:0] _RAND_4235;
  reg [31:0] _RAND_4236;
  reg [31:0] _RAND_4237;
  reg [31:0] _RAND_4238;
  reg [31:0] _RAND_4239;
  reg [31:0] _RAND_4240;
  reg [31:0] _RAND_4241;
  reg [31:0] _RAND_4242;
  reg [31:0] _RAND_4243;
  reg [31:0] _RAND_4244;
  reg [31:0] _RAND_4245;
  reg [31:0] _RAND_4246;
  reg [31:0] _RAND_4247;
  reg [31:0] _RAND_4248;
  reg [31:0] _RAND_4249;
  reg [31:0] _RAND_4250;
  reg [31:0] _RAND_4251;
  reg [31:0] _RAND_4252;
  reg [31:0] _RAND_4253;
  reg [31:0] _RAND_4254;
  reg [31:0] _RAND_4255;
  reg [31:0] _RAND_4256;
  reg [31:0] _RAND_4257;
  reg [31:0] _RAND_4258;
  reg [31:0] _RAND_4259;
  reg [31:0] _RAND_4260;
  reg [31:0] _RAND_4261;
  reg [31:0] _RAND_4262;
  reg [31:0] _RAND_4263;
  reg [31:0] _RAND_4264;
  reg [31:0] _RAND_4265;
  reg [31:0] _RAND_4266;
  reg [31:0] _RAND_4267;
  reg [31:0] _RAND_4268;
  reg [31:0] _RAND_4269;
  reg [31:0] _RAND_4270;
  reg [31:0] _RAND_4271;
  reg [31:0] _RAND_4272;
  reg [31:0] _RAND_4273;
  reg [31:0] _RAND_4274;
  reg [31:0] _RAND_4275;
  reg [31:0] _RAND_4276;
  reg [31:0] _RAND_4277;
  reg [31:0] _RAND_4278;
  reg [31:0] _RAND_4279;
  reg [31:0] _RAND_4280;
  reg [31:0] _RAND_4281;
  reg [31:0] _RAND_4282;
  reg [31:0] _RAND_4283;
  reg [31:0] _RAND_4284;
  reg [31:0] _RAND_4285;
  reg [31:0] _RAND_4286;
  reg [31:0] _RAND_4287;
  reg [31:0] _RAND_4288;
  reg [31:0] _RAND_4289;
  reg [31:0] _RAND_4290;
  reg [31:0] _RAND_4291;
  reg [31:0] _RAND_4292;
  reg [31:0] _RAND_4293;
  reg [31:0] _RAND_4294;
  reg [31:0] _RAND_4295;
  reg [31:0] _RAND_4296;
  reg [31:0] _RAND_4297;
  reg [31:0] _RAND_4298;
  reg [31:0] _RAND_4299;
  reg [31:0] _RAND_4300;
  reg [31:0] _RAND_4301;
  reg [31:0] _RAND_4302;
  reg [31:0] _RAND_4303;
  reg [31:0] _RAND_4304;
  reg [31:0] _RAND_4305;
  reg [31:0] _RAND_4306;
  reg [31:0] _RAND_4307;
  reg [31:0] _RAND_4308;
  reg [31:0] _RAND_4309;
  reg [31:0] _RAND_4310;
  reg [31:0] _RAND_4311;
  reg [31:0] _RAND_4312;
  reg [31:0] _RAND_4313;
  reg [31:0] _RAND_4314;
  reg [31:0] _RAND_4315;
  reg [31:0] _RAND_4316;
  reg [31:0] _RAND_4317;
  reg [31:0] _RAND_4318;
  reg [31:0] _RAND_4319;
  reg [31:0] _RAND_4320;
  reg [31:0] _RAND_4321;
  reg [31:0] _RAND_4322;
  reg [31:0] _RAND_4323;
  reg [31:0] _RAND_4324;
  reg [31:0] _RAND_4325;
  reg [31:0] _RAND_4326;
  reg [31:0] _RAND_4327;
  reg [31:0] _RAND_4328;
  reg [31:0] _RAND_4329;
  reg [31:0] _RAND_4330;
  reg [31:0] _RAND_4331;
  reg [31:0] _RAND_4332;
  reg [31:0] _RAND_4333;
  reg [31:0] _RAND_4334;
  reg [31:0] _RAND_4335;
  reg [31:0] _RAND_4336;
  reg [31:0] _RAND_4337;
  reg [31:0] _RAND_4338;
  reg [31:0] _RAND_4339;
  reg [31:0] _RAND_4340;
  reg [31:0] _RAND_4341;
  reg [31:0] _RAND_4342;
  reg [31:0] _RAND_4343;
  reg [31:0] _RAND_4344;
  reg [31:0] _RAND_4345;
  reg [31:0] _RAND_4346;
  reg [31:0] _RAND_4347;
  reg [31:0] _RAND_4348;
  reg [31:0] _RAND_4349;
  reg [31:0] _RAND_4350;
  reg [31:0] _RAND_4351;
  reg [31:0] _RAND_4352;
  reg [31:0] _RAND_4353;
  reg [31:0] _RAND_4354;
  reg [31:0] _RAND_4355;
  reg [31:0] _RAND_4356;
  reg [31:0] _RAND_4357;
  reg [31:0] _RAND_4358;
  reg [31:0] _RAND_4359;
  reg [31:0] _RAND_4360;
  reg [31:0] _RAND_4361;
  reg [31:0] _RAND_4362;
  reg [31:0] _RAND_4363;
  reg [31:0] _RAND_4364;
  reg [31:0] _RAND_4365;
  reg [31:0] _RAND_4366;
  reg [31:0] _RAND_4367;
  reg [31:0] _RAND_4368;
  reg [31:0] _RAND_4369;
  reg [31:0] _RAND_4370;
  reg [31:0] _RAND_4371;
  reg [31:0] _RAND_4372;
  reg [31:0] _RAND_4373;
  reg [31:0] _RAND_4374;
  reg [31:0] _RAND_4375;
  reg [31:0] _RAND_4376;
  reg [31:0] _RAND_4377;
  reg [31:0] _RAND_4378;
  reg [31:0] _RAND_4379;
  reg [31:0] _RAND_4380;
  reg [31:0] _RAND_4381;
  reg [31:0] _RAND_4382;
  reg [31:0] _RAND_4383;
  reg [31:0] _RAND_4384;
  reg [31:0] _RAND_4385;
  reg [31:0] _RAND_4386;
  reg [31:0] _RAND_4387;
  reg [31:0] _RAND_4388;
  reg [31:0] _RAND_4389;
  reg [31:0] _RAND_4390;
  reg [31:0] _RAND_4391;
  reg [31:0] _RAND_4392;
  reg [31:0] _RAND_4393;
  reg [31:0] _RAND_4394;
  reg [31:0] _RAND_4395;
  reg [31:0] _RAND_4396;
  reg [31:0] _RAND_4397;
  reg [31:0] _RAND_4398;
  reg [31:0] _RAND_4399;
  reg [31:0] _RAND_4400;
  reg [31:0] _RAND_4401;
  reg [31:0] _RAND_4402;
  reg [31:0] _RAND_4403;
  reg [31:0] _RAND_4404;
  reg [31:0] _RAND_4405;
  reg [31:0] _RAND_4406;
  reg [31:0] _RAND_4407;
  reg [31:0] _RAND_4408;
  reg [31:0] _RAND_4409;
  reg [31:0] _RAND_4410;
  reg [31:0] _RAND_4411;
  reg [31:0] _RAND_4412;
  reg [31:0] _RAND_4413;
  reg [31:0] _RAND_4414;
  reg [31:0] _RAND_4415;
  reg [31:0] _RAND_4416;
  reg [31:0] _RAND_4417;
  reg [31:0] _RAND_4418;
  reg [31:0] _RAND_4419;
  reg [31:0] _RAND_4420;
  reg [31:0] _RAND_4421;
  reg [31:0] _RAND_4422;
  reg [31:0] _RAND_4423;
  reg [31:0] _RAND_4424;
  reg [31:0] _RAND_4425;
  reg [31:0] _RAND_4426;
  reg [31:0] _RAND_4427;
  reg [31:0] _RAND_4428;
  reg [31:0] _RAND_4429;
  reg [31:0] _RAND_4430;
  reg [31:0] _RAND_4431;
  reg [31:0] _RAND_4432;
  reg [31:0] _RAND_4433;
  reg [31:0] _RAND_4434;
  reg [31:0] _RAND_4435;
  reg [31:0] _RAND_4436;
  reg [31:0] _RAND_4437;
  reg [31:0] _RAND_4438;
  reg [31:0] _RAND_4439;
  reg [31:0] _RAND_4440;
  reg [31:0] _RAND_4441;
  reg [31:0] _RAND_4442;
  reg [31:0] _RAND_4443;
  reg [31:0] _RAND_4444;
  reg [31:0] _RAND_4445;
  reg [31:0] _RAND_4446;
  reg [31:0] _RAND_4447;
  reg [31:0] _RAND_4448;
  reg [31:0] _RAND_4449;
  reg [31:0] _RAND_4450;
  reg [31:0] _RAND_4451;
  reg [31:0] _RAND_4452;
  reg [31:0] _RAND_4453;
  reg [31:0] _RAND_4454;
  reg [31:0] _RAND_4455;
  reg [31:0] _RAND_4456;
  reg [31:0] _RAND_4457;
  reg [31:0] _RAND_4458;
  reg [31:0] _RAND_4459;
  reg [31:0] _RAND_4460;
  reg [31:0] _RAND_4461;
  reg [31:0] _RAND_4462;
  reg [31:0] _RAND_4463;
  reg [31:0] _RAND_4464;
  reg [31:0] _RAND_4465;
  reg [31:0] _RAND_4466;
  reg [31:0] _RAND_4467;
  reg [31:0] _RAND_4468;
  reg [31:0] _RAND_4469;
  reg [31:0] _RAND_4470;
  reg [31:0] _RAND_4471;
  reg [31:0] _RAND_4472;
  reg [31:0] _RAND_4473;
  reg [31:0] _RAND_4474;
  reg [31:0] _RAND_4475;
  reg [31:0] _RAND_4476;
  reg [31:0] _RAND_4477;
  reg [31:0] _RAND_4478;
  reg [31:0] _RAND_4479;
  reg [31:0] _RAND_4480;
  reg [31:0] _RAND_4481;
  reg [31:0] _RAND_4482;
  reg [31:0] _RAND_4483;
  reg [31:0] _RAND_4484;
  reg [31:0] _RAND_4485;
  reg [31:0] _RAND_4486;
  reg [31:0] _RAND_4487;
  reg [31:0] _RAND_4488;
  reg [31:0] _RAND_4489;
  reg [31:0] _RAND_4490;
  reg [31:0] _RAND_4491;
  reg [31:0] _RAND_4492;
  reg [31:0] _RAND_4493;
  reg [31:0] _RAND_4494;
  reg [31:0] _RAND_4495;
  reg [31:0] _RAND_4496;
  reg [31:0] _RAND_4497;
  reg [31:0] _RAND_4498;
  reg [31:0] _RAND_4499;
  reg [31:0] _RAND_4500;
  reg [31:0] _RAND_4501;
  reg [31:0] _RAND_4502;
  reg [31:0] _RAND_4503;
  reg [31:0] _RAND_4504;
  reg [31:0] _RAND_4505;
  reg [31:0] _RAND_4506;
  reg [31:0] _RAND_4507;
  reg [31:0] _RAND_4508;
  reg [31:0] _RAND_4509;
  reg [31:0] _RAND_4510;
  reg [31:0] _RAND_4511;
  reg [31:0] _RAND_4512;
  reg [31:0] _RAND_4513;
  reg [31:0] _RAND_4514;
  reg [31:0] _RAND_4515;
  reg [31:0] _RAND_4516;
  reg [31:0] _RAND_4517;
  reg [31:0] _RAND_4518;
  reg [31:0] _RAND_4519;
  reg [31:0] _RAND_4520;
  reg [31:0] _RAND_4521;
  reg [31:0] _RAND_4522;
  reg [31:0] _RAND_4523;
  reg [31:0] _RAND_4524;
  reg [31:0] _RAND_4525;
  reg [31:0] _RAND_4526;
  reg [31:0] _RAND_4527;
  reg [31:0] _RAND_4528;
  reg [31:0] _RAND_4529;
  reg [31:0] _RAND_4530;
  reg [31:0] _RAND_4531;
  reg [31:0] _RAND_4532;
  reg [31:0] _RAND_4533;
  reg [31:0] _RAND_4534;
  reg [31:0] _RAND_4535;
  reg [31:0] _RAND_4536;
  reg [31:0] _RAND_4537;
  reg [31:0] _RAND_4538;
  reg [31:0] _RAND_4539;
  reg [31:0] _RAND_4540;
  reg [31:0] _RAND_4541;
  reg [31:0] _RAND_4542;
  reg [31:0] _RAND_4543;
  reg [31:0] _RAND_4544;
  reg [31:0] _RAND_4545;
  reg [31:0] _RAND_4546;
  reg [31:0] _RAND_4547;
  reg [31:0] _RAND_4548;
  reg [31:0] _RAND_4549;
  reg [31:0] _RAND_4550;
  reg [31:0] _RAND_4551;
  reg [31:0] _RAND_4552;
  reg [31:0] _RAND_4553;
  reg [31:0] _RAND_4554;
  reg [31:0] _RAND_4555;
  reg [31:0] _RAND_4556;
  reg [31:0] _RAND_4557;
  reg [31:0] _RAND_4558;
  reg [31:0] _RAND_4559;
  reg [31:0] _RAND_4560;
  reg [31:0] _RAND_4561;
  reg [31:0] _RAND_4562;
  reg [31:0] _RAND_4563;
  reg [31:0] _RAND_4564;
  reg [31:0] _RAND_4565;
  reg [31:0] _RAND_4566;
  reg [31:0] _RAND_4567;
  reg [31:0] _RAND_4568;
  reg [31:0] _RAND_4569;
  reg [31:0] _RAND_4570;
  reg [31:0] _RAND_4571;
  reg [31:0] _RAND_4572;
  reg [31:0] _RAND_4573;
  reg [31:0] _RAND_4574;
  reg [31:0] _RAND_4575;
  reg [31:0] _RAND_4576;
  reg [31:0] _RAND_4577;
  reg [31:0] _RAND_4578;
  reg [31:0] _RAND_4579;
  reg [31:0] _RAND_4580;
  reg [31:0] _RAND_4581;
  reg [31:0] _RAND_4582;
  reg [31:0] _RAND_4583;
  reg [31:0] _RAND_4584;
  reg [31:0] _RAND_4585;
  reg [31:0] _RAND_4586;
  reg [31:0] _RAND_4587;
  reg [31:0] _RAND_4588;
  reg [31:0] _RAND_4589;
  reg [31:0] _RAND_4590;
  reg [31:0] _RAND_4591;
  reg [31:0] _RAND_4592;
  reg [31:0] _RAND_4593;
  reg [31:0] _RAND_4594;
  reg [31:0] _RAND_4595;
  reg [31:0] _RAND_4596;
  reg [31:0] _RAND_4597;
  reg [31:0] _RAND_4598;
  reg [31:0] _RAND_4599;
  reg [31:0] _RAND_4600;
  reg [31:0] _RAND_4601;
  reg [31:0] _RAND_4602;
  reg [31:0] _RAND_4603;
  reg [31:0] _RAND_4604;
  reg [31:0] _RAND_4605;
  reg [31:0] _RAND_4606;
  reg [31:0] _RAND_4607;
`endif // RANDOMIZE_REG_INIT
  wire  mesh_0_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_0_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_0_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_0_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_0_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_0_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_1_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_1_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_1_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_1_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_1_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_2_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_2_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_2_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_2_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_2_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_3_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_3_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_3_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_3_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_3_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_4_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_4_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_4_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_4_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_4_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_5_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_5_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_5_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_5_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_5_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_6_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_6_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_6_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_6_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_6_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_7_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_7_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_7_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_7_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_7_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_8_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_8_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_8_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_8_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_8_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_9_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_9_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_9_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_9_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_9_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_10_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_10_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_10_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_10_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_10_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_11_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_11_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_11_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_11_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_11_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_12_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_12_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_12_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_12_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_12_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_13_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_13_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_13_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_13_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_13_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_14_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_14_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_14_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_14_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_14_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_0_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_0_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_0_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_0_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_0_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_0_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_1_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_1_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_1_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_1_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_1_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_1_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_2_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_2_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_2_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_2_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_2_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_2_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_3_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_3_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_3_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_3_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_3_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_3_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_4_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_4_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_4_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_4_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_4_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_4_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_5_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_5_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_5_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_5_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_5_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_5_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_6_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_6_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_6_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_6_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_6_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_6_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_7_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_7_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_7_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_7_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_7_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_7_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_8_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_8_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_8_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_8_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_8_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_8_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_9_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_9_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_9_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_9_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_9_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_9_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_10_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_10_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_10_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_10_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_10_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_10_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_11_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_11_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_11_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_11_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_11_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_11_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_12_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_12_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_12_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_12_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_12_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_12_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_13_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_13_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_13_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_13_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_13_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_13_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_14_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_14_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_14_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_14_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_14_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_14_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_clock; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_15_io_in_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_15_io_in_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_in_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_in_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_in_d_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_in_d_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_15_io_in_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_15_io_in_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_15_io_in_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_15_io_in_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_15_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [7:0] mesh_15_15_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [19:0] mesh_15_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [4:0] mesh_15_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire [1:0] mesh_15_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_in_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  wire  mesh_15_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 39:71]
  reg [7:0] r__0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r__1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_1_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_1_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_2_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_2_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_3_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_3_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_4_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_4_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_5_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_5_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_6_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_6_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_7_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_7_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_8_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_8_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_9_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_9_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_10_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_10_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_11_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_11_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_12_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_12_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_13_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_13_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_14_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_14_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_15_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_15_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_16_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_16_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_17_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_17_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_18_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_18_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_19_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_19_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_20_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_20_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_21_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_21_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_22_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_22_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_23_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_23_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_24_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_24_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_25_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_25_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_26_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_26_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_27_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_27_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_28_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_28_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_29_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_29_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_30_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_30_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_31_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_31_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_32_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_32_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_33_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_33_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_34_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_34_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_35_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_35_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_36_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_36_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_37_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_37_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_38_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_38_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_39_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_39_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_40_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_40_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_41_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_41_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_42_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_42_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_43_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_43_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_44_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_44_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_45_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_45_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_46_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_46_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_47_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_47_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_48_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_48_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_49_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_49_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_50_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_50_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_51_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_51_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_52_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_52_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_53_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_53_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_54_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_54_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_55_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_55_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_56_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_56_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_57_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_57_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_58_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_58_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_59_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_59_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_60_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_60_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_61_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_61_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_62_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_62_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_63_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_63_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_64_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_64_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_65_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_65_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_66_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_66_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_67_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_67_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_68_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_68_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_69_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_69_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_70_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_70_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_71_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_71_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_72_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_72_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_73_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_73_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_74_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_74_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_75_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_75_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_76_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_76_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_77_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_77_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_78_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_78_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_79_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_79_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_80_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_80_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_81_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_81_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_82_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_82_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_83_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_83_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_84_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_84_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_85_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_85_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_86_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_86_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_87_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_87_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_88_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_88_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_89_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_89_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_90_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_90_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_91_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_91_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_92_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_92_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_93_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_93_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_94_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_94_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_95_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_95_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_96_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_96_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_97_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_97_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_98_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_98_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_99_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_99_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_100_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_100_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_101_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_101_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_102_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_102_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_103_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_103_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_104_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_104_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_105_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_105_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_106_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_106_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_107_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_107_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_108_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_108_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_109_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_109_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_110_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_110_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_111_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_111_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_112_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_112_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_113_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_113_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_114_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_114_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_115_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_115_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_116_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_116_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_117_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_117_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_118_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_118_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_119_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_119_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_120_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_120_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_121_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_121_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_122_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_122_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_123_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_123_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_124_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_124_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_125_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_125_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_126_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_126_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_127_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_127_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_128_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_128_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_129_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_129_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_130_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_130_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_131_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_131_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_132_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_132_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_133_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_133_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_134_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_134_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_135_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_135_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_136_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_136_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_137_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_137_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_138_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_138_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_139_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_139_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_140_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_140_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_141_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_141_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_142_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_142_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_143_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_143_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_144_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_144_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_145_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_145_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_146_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_146_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_147_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_147_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_148_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_148_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_149_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_149_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_150_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_150_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_151_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_151_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_152_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_152_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_153_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_153_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_154_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_154_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_155_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_155_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_156_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_156_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_157_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_157_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_158_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_158_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_159_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_159_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_160_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_160_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_161_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_161_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_162_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_162_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_163_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_163_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_164_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_164_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_165_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_165_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_166_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_166_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_167_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_167_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_168_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_168_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_169_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_169_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_170_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_170_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_171_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_171_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_172_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_172_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_173_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_173_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_174_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_174_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_175_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_175_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_176_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_176_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_177_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_177_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_178_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_178_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_179_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_179_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_180_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_180_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_181_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_181_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_182_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_182_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_183_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_183_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_184_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_184_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_185_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_185_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_186_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_186_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_187_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_187_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_188_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_188_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_189_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_189_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_190_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_190_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_191_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_191_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_192_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_192_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_193_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_193_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_194_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_194_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_195_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_195_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_196_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_196_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_197_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_197_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_198_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_198_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_199_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_199_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_200_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_200_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_201_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_201_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_202_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_202_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_203_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_203_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_204_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_204_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_205_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_205_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_206_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_206_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_207_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_207_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_208_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_208_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_209_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_209_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_210_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_210_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_211_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_211_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_212_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_212_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_213_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_213_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_214_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_214_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_215_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_215_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_216_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_216_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_217_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_217_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_218_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_218_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_219_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_219_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_220_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_220_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_221_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_221_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_222_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_222_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_223_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_223_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_224_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_224_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_225_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_225_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_226_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_226_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_227_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_227_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_228_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_228_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_229_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_229_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_230_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_230_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_231_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_231_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_232_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_232_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_233_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_233_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_234_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_234_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_235_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_235_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_236_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_236_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_237_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_237_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_238_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_238_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_239_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_239_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_240_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_240_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_241_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_241_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_242_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_242_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_243_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_243_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_244_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_244_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_245_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_245_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_246_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_246_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_247_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_247_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_248_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_248_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_249_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_249_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_250_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_250_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_251_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_251_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_252_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_252_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_253_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_253_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_254_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_254_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_255_0; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] r_255_1; // @[src/main/scala/gemmini/Mesh.scala 53:38]
  reg [7:0] pipe_b__0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b__1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_1_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_1_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_2_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_2_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_3_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_3_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_4_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_4_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_5_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_5_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_6_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_6_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_7_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_7_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_8_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_8_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_9_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_9_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_10_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_10_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_11_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_11_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_12_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_12_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_13_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_13_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_14_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_14_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_15_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_15_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_16_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_16_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_17_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_17_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_18_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_18_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_19_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_19_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_20_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_20_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_21_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_21_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_22_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_22_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_23_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_23_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_24_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_24_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_25_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_25_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_26_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_26_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_27_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_27_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_28_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_28_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_29_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_29_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_30_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_30_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_31_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_31_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_32_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_32_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_33_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_33_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_34_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_34_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_35_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_35_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_36_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_36_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_37_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_37_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_38_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_38_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_39_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_39_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_40_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_40_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_41_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_41_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_42_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_42_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_43_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_43_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_44_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_44_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_45_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_45_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_46_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_46_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_47_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_47_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_48_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_48_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_49_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_49_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_50_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_50_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_51_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_51_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_52_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_52_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_53_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_53_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_54_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_54_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_55_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_55_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_56_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_56_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_57_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_57_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_58_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_58_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_59_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_59_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_60_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_60_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_61_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_61_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_62_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_62_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_63_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_63_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_64_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_64_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_65_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_65_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_66_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_66_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_67_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_67_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_68_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_68_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_69_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_69_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_70_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_70_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_71_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_71_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_72_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_72_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_73_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_73_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_74_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_74_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_75_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_75_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_76_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_76_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_77_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_77_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_78_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_78_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_79_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_79_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_80_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_80_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_81_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_81_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_82_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_82_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_83_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_83_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_84_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_84_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_85_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_85_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_86_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_86_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_87_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_87_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_88_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_88_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_89_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_89_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_90_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_90_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_91_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_91_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_92_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_92_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_93_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_93_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_94_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_94_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_95_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_95_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_96_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_96_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_97_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_97_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_98_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_98_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_99_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_99_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_100_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_100_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_101_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_101_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_102_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_102_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_103_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_103_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_104_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_104_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_105_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_105_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_106_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_106_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_107_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_107_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_108_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_108_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_109_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_109_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_110_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_110_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_111_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_111_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_112_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_112_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_113_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_113_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_114_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_114_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_115_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_115_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_116_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_116_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_117_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_117_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_118_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_118_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_119_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_119_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_120_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_120_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_121_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_121_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_122_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_122_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_123_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_123_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_124_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_124_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_125_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_125_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_126_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_126_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_127_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_127_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_128_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_128_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_129_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_129_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_130_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_130_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_131_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_131_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_132_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_132_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_133_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_133_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_134_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_134_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_135_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_135_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_136_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_136_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_137_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_137_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_138_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_138_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_139_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_139_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_140_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_140_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_141_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_141_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_142_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_142_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_143_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_143_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_144_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_144_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_145_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_145_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_146_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_146_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_147_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_147_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_148_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_148_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_149_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_149_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_150_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_150_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_151_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_151_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_152_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_152_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_153_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_153_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_154_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_154_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_155_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_155_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_156_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_156_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_157_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_157_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_158_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_158_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_159_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_159_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_160_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_160_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_161_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_161_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_162_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_162_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_163_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_163_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_164_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_164_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_165_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_165_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_166_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_166_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_167_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_167_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_168_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_168_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_169_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_169_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_170_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_170_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_171_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_171_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_172_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_172_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_173_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_173_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_174_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_174_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_175_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_175_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_176_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_176_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_177_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_177_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_178_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_178_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_179_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_179_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_180_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_180_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_181_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_181_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_182_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_182_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_183_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_183_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_184_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_184_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_185_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_185_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_186_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_186_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_187_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_187_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_188_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_188_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_189_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_189_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_190_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_190_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_191_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_191_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_192_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_192_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_193_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_193_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_194_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_194_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_195_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_195_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_196_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_196_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_197_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_197_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_198_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_198_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_199_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_199_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_200_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_200_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_201_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_201_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_202_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_202_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_203_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_203_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_204_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_204_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_205_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_205_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_206_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_206_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_207_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_207_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_208_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_208_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_209_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_209_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_210_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_210_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_211_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_211_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_212_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_212_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_213_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_213_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_214_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_214_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_215_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_215_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_216_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_216_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_217_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_217_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_218_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_218_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_219_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_219_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_220_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_220_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_221_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_221_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_222_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_222_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_223_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_223_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_224_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_224_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_225_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_225_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_226_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_226_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_227_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_227_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_228_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_228_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_229_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_229_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_230_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_230_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_231_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_231_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_232_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_232_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_233_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_233_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_234_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_234_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_235_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_235_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_236_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_236_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_237_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_237_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_238_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_238_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_239_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_239_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_240_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_240_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_241_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_241_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_242_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_242_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_243_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_243_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_244_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_244_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_245_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_245_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_246_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_246_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_247_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_247_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_248_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_248_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_249_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_249_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_250_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_250_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_251_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_251_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_252_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_252_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_253_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_253_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_254_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_254_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_255_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_255_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_256_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_256_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_257_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_257_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_258_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_258_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_259_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_259_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_260_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_260_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_261_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_261_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_262_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_262_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_263_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_263_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_264_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_264_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_265_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_265_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_266_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_266_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_267_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_267_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_268_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_268_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_269_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_269_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_270_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_270_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_271_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_271_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_272_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_272_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_273_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_273_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_274_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_274_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_275_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_275_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_276_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_276_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_277_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_277_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_278_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_278_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_279_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_279_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_280_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_280_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_281_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_281_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_282_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_282_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_283_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_283_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_284_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_284_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_285_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_285_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_286_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_286_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_287_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_287_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_288_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_288_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_289_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_289_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_290_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_290_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_291_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_291_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_292_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_292_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_293_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_293_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_294_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_294_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_295_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_295_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_296_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_296_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_297_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_297_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_298_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_298_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_299_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_299_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_300_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_300_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_301_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_301_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_302_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_302_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_303_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_303_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_304_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_304_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_305_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_305_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_306_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_306_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_307_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_307_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_308_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_308_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_309_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_309_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_310_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_310_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_311_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_311_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_312_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_312_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_313_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_313_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_314_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_314_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_315_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_315_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_316_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_316_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_317_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_317_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_318_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_318_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_319_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_319_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_320_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_320_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_321_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_321_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_322_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_322_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_323_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_323_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_324_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_324_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_325_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_325_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_326_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_326_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_327_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_327_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_328_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_328_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_329_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_329_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_330_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_330_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_331_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_331_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_332_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_332_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_333_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_333_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_334_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_334_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_335_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_335_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_336_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_336_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_337_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_337_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_338_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_338_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_339_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_339_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_340_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_340_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_341_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_341_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_342_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_342_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_343_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_343_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_344_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_344_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_345_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_345_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_346_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_346_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_347_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_347_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_348_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_348_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_349_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_349_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_350_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_350_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_351_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_351_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_352_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_352_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_353_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_353_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_354_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_354_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_355_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_355_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_356_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_356_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_357_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_357_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_358_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_358_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_359_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_359_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_360_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_360_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_361_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_361_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_362_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_362_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_363_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_363_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_364_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_364_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_365_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_365_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_366_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_366_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_367_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_367_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_368_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_368_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_369_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_369_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_370_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_370_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_371_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_371_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_372_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_372_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_373_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_373_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_374_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_374_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_375_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_375_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_376_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_376_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_377_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_377_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_378_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_378_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_379_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_379_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_380_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_380_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_381_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_381_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_382_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_382_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_383_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_383_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_384_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_384_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_385_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_385_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_386_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_386_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_387_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_387_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_388_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_388_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_389_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_389_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_390_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_390_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_391_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_391_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_392_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_392_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_393_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_393_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_394_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_394_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_395_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_395_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_396_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_396_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_397_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_397_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_398_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_398_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_399_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_399_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_400_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_400_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_401_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_401_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_402_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_402_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_403_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_403_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_404_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_404_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_405_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_405_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_406_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_406_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_407_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_407_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_408_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_408_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_409_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_409_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_410_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_410_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_411_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_411_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_412_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_412_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_413_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_413_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_414_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_414_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_415_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_415_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_416_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_416_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_417_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_417_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_418_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_418_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_419_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_419_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_420_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_420_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_421_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_421_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_422_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_422_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_423_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_423_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_424_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_424_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_425_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_425_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_426_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_426_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_427_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_427_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_428_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_428_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_429_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_429_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_430_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_430_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_431_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_431_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_432_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_432_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_433_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_433_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_434_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_434_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_435_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_435_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_436_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_436_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_437_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_437_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_438_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_438_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_439_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_439_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_440_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_440_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_441_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_441_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_442_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_442_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_443_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_443_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_444_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_444_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_445_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_445_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_446_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_446_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_447_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_447_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_448_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_448_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_449_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_449_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_450_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_450_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_451_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_451_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_452_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_452_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_453_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_453_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_454_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_454_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_455_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_455_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_456_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_456_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_457_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_457_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_458_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_458_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_459_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_459_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_460_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_460_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_461_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_461_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_462_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_462_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_463_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_463_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_464_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_464_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_465_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_465_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_466_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_466_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_467_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_467_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_468_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_468_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_469_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_469_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_470_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_470_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_471_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_471_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_472_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_472_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_473_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_473_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_474_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_474_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_475_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_475_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_476_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_476_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_477_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_477_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_478_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_478_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_479_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_479_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_480_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_480_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_481_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_481_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_482_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_482_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_483_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_483_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_484_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_484_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_485_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_485_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_486_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_486_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_487_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_487_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_488_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_488_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_489_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_489_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_490_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_490_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_491_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_491_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_492_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_492_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_493_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_493_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_494_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_494_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_495_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_495_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_496_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [7:0] pipe_b_496_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_497_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_497_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_498_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_498_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_499_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_499_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_500_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_500_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_501_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_501_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_502_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_502_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_503_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_503_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_504_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_504_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_505_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_505_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_506_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_506_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_507_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_507_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_508_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_508_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_509_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_509_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_510_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_510_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_511_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [19:0] pipe_b_511_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_0_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_0_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_1_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_1_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_2_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_2_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_3_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_3_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_4_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_4_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_5_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_5_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_6_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_6_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_7_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_7_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_8_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_8_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_9_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_9_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_10_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_10_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_11_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_11_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_12_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_12_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_13_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_13_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_14_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_14_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg [4:0] mesh_15_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  mesh_15_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
  reg  r_256_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_256_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_257_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_257_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_258_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_258_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_259_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_259_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_260_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_260_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_261_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_261_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_262_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_262_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_263_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_263_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_264_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_264_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_265_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_265_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_266_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_266_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_267_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_267_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_268_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_268_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_269_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_269_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_270_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_270_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_271_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_271_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_272_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_272_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_273_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_273_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_274_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_274_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_275_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_275_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_276_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_276_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_277_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_277_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_278_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_278_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_279_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_279_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_280_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_280_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_281_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_281_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_282_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_282_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_283_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_283_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_284_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_284_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_285_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_285_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_286_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_286_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_287_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_287_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_288_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_288_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_289_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_289_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_290_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_290_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_291_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_291_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_292_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_292_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_293_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_293_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_294_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_294_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_295_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_295_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_296_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_296_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_297_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_297_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_298_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_298_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_299_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_299_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_300_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_300_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_301_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_301_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_302_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_302_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_303_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_303_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_304_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_304_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_305_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_305_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_306_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_306_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_307_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_307_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_308_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_308_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_309_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_309_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_310_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_310_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_311_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_311_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_312_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_312_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_313_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_313_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_314_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_314_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_315_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_315_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_316_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_316_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_317_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_317_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_318_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_318_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_319_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_319_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_320_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_320_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_321_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_321_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_322_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_322_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_323_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_323_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_324_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_324_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_325_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_325_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_326_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_326_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_327_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_327_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_328_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_328_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_329_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_329_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_330_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_330_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_331_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_331_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_332_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_332_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_333_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_333_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_334_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_334_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_335_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_335_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_336_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_336_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_337_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_337_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_338_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_338_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_339_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_339_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_340_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_340_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_341_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_341_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_342_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_342_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_343_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_343_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_344_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_344_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_345_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_345_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_346_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_346_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_347_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_347_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_348_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_348_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_349_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_349_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_350_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_350_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_351_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_351_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_352_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_352_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_353_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_353_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_354_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_354_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_355_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_355_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_356_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_356_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_357_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_357_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_358_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_358_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_359_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_359_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_360_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_360_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_361_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_361_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_362_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_362_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_363_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_363_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_364_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_364_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_365_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_365_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_366_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_366_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_367_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_367_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_368_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_368_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_369_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_369_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_370_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_370_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_371_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_371_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_372_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_372_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_373_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_373_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_374_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_374_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_375_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_375_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_376_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_376_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_377_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_377_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_378_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_378_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_379_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_379_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_380_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_380_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_381_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_381_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_382_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_382_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_383_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_383_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_384_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_384_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_385_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_385_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_386_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_386_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_387_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_387_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_388_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_388_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_389_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_389_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_390_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_390_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_391_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_391_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_392_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_392_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_393_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_393_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_394_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_394_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_395_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_395_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_396_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_396_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_397_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_397_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_398_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_398_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_399_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_399_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_400_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_400_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_401_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_401_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_402_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_402_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_403_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_403_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_404_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_404_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_405_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_405_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_406_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_406_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_407_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_407_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_408_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_408_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_409_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_409_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_410_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_410_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_411_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_411_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_412_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_412_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_413_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_413_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_414_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_414_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_415_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_415_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_416_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_416_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_417_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_417_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_418_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_418_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_419_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_419_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_420_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_420_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_421_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_421_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_422_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_422_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_423_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_423_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_424_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_424_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_425_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_425_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_426_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_426_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_427_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_427_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_428_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_428_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_429_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_429_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_430_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_430_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_431_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_431_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_432_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_432_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_433_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_433_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_434_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_434_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_435_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_435_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_436_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_436_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_437_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_437_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_438_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_438_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_439_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_439_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_440_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_440_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_441_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_441_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_442_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_442_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_443_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_443_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_444_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_444_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_445_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_445_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_446_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_446_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_447_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_447_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_448_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_448_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_449_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_449_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_450_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_450_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_451_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_451_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_452_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_452_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_453_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_453_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_454_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_454_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_455_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_455_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_456_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_456_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_457_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_457_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_458_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_458_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_459_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_459_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_460_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_460_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_461_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_461_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_462_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_462_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_463_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_463_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_464_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_464_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_465_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_465_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_466_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_466_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_467_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_467_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_468_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_468_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_469_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_469_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_470_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_470_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_471_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_471_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_472_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_472_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_473_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_473_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_474_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_474_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_475_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_475_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_476_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_476_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_477_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_477_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_478_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_478_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_479_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_479_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_480_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_480_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_481_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_481_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_482_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_482_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_483_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_483_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_484_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_484_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_485_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_485_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_486_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_486_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_487_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_487_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_488_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_488_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_489_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_489_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_490_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_490_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_491_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_491_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_492_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_492_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_493_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_493_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_494_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_494_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_495_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_495_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_496_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_496_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_497_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_497_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_498_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_498_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_499_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_499_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_500_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_500_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_501_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_501_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_502_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_502_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_503_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_503_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_504_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_504_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_505_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_505_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_506_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_506_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_507_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_507_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_508_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_508_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_509_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_509_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_510_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_510_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_511_0; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg  r_511_1; // @[src/main/scala/gemmini/Mesh.scala 94:42]
  reg [1:0] r_512_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_512_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_513_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_513_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_514_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_514_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_515_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_515_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_516_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_516_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_517_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_517_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_518_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_518_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_519_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_519_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_520_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_520_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_521_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_521_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_522_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_522_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_523_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_523_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_524_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_524_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_525_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_525_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_526_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_526_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_527_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_527_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_528_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_528_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_529_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_529_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_530_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_530_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_531_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_531_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_532_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_532_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_533_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_533_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_534_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_534_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_535_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_535_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_536_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_536_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_537_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_537_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_538_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_538_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_539_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_539_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_540_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_540_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_541_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_541_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_542_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_542_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_543_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_543_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_544_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_544_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_545_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_545_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_546_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_546_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_547_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_547_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_548_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_548_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_549_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_549_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_550_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_550_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_551_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_551_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_552_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_552_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_553_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_553_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_554_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_554_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_555_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_555_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_556_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_556_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_557_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_557_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_558_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_558_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_559_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_559_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_560_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_560_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_561_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_561_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_562_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_562_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_563_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_563_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_564_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_564_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_565_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_565_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_566_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_566_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_567_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_567_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_568_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_568_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_569_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_569_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_570_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_570_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_571_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_571_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_572_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_572_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_573_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_573_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_574_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_574_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_575_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_575_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_576_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_576_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_577_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_577_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_578_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_578_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_579_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_579_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_580_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_580_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_581_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_581_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_582_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_582_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_583_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_583_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_584_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_584_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_585_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_585_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_586_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_586_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_587_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_587_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_588_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_588_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_589_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_589_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_590_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_590_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_591_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_591_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_592_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_592_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_593_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_593_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_594_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_594_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_595_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_595_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_596_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_596_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_597_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_597_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_598_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_598_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_599_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_599_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_600_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_600_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_601_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_601_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_602_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_602_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_603_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_603_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_604_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_604_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_605_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_605_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_606_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_606_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_607_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_607_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_608_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_608_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_609_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_609_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_610_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_610_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_611_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_611_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_612_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_612_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_613_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_613_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_614_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_614_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_615_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_615_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_616_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_616_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_617_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_617_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_618_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_618_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_619_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_619_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_620_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_620_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_621_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_621_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_622_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_622_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_623_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_623_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_624_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_624_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_625_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_625_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_626_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_626_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_627_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_627_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_628_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_628_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_629_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_629_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_630_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_630_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_631_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_631_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_632_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_632_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_633_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_633_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_634_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_634_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_635_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_635_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_636_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_636_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_637_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_637_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_638_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_638_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_639_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_639_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_640_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_640_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_641_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_641_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_642_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_642_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_643_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_643_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_644_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_644_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_645_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_645_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_646_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_646_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_647_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_647_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_648_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_648_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_649_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_649_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_650_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_650_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_651_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_651_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_652_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_652_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_653_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_653_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_654_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_654_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_655_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_655_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_656_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_656_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_657_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_657_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_658_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_658_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_659_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_659_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_660_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_660_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_661_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_661_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_662_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_662_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_663_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_663_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_664_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_664_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_665_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_665_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_666_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_666_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_667_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_667_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_668_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_668_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_669_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_669_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_670_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_670_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_671_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_671_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_672_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_672_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_673_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_673_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_674_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_674_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_675_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_675_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_676_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_676_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_677_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_677_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_678_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_678_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_679_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_679_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_680_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_680_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_681_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_681_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_682_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_682_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_683_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_683_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_684_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_684_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_685_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_685_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_686_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_686_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_687_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_687_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_688_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_688_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_689_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_689_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_690_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_690_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_691_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_691_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_692_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_692_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_693_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_693_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_694_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_694_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_695_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_695_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_696_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_696_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_697_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_697_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_698_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_698_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_699_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_699_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_700_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_700_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_701_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_701_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_702_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_702_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_703_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_703_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_704_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_704_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_705_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_705_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_706_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_706_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_707_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_707_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_708_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_708_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_709_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_709_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_710_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_710_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_711_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_711_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_712_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_712_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_713_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_713_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_714_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_714_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_715_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_715_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_716_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_716_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_717_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_717_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_718_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_718_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_719_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_719_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_720_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_720_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_721_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_721_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_722_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_722_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_723_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_723_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_724_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_724_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_725_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_725_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_726_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_726_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_727_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_727_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_728_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_728_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_729_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_729_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_730_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_730_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_731_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_731_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_732_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_732_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_733_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_733_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_734_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_734_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_735_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_735_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_736_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_736_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_737_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_737_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_738_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_738_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_739_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_739_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_740_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_740_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_741_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_741_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_742_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_742_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_743_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_743_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_744_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_744_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_745_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_745_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_746_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_746_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_747_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_747_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_748_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_748_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_749_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_749_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_750_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_750_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_751_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_751_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_752_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_752_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_753_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_753_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_754_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_754_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_755_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_755_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_756_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_756_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_757_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_757_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_758_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_758_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_759_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_759_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_760_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_760_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_761_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_761_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_762_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_762_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_763_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_763_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_764_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_764_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_765_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_765_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_766_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_766_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_767_0; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg [1:0] r_767_1; // @[src/main/scala/gemmini/Mesh.scala 103:39]
  reg  r_768_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_768_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_769_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_769_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_770_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_770_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_771_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_771_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_772_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_772_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_773_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_773_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_774_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_774_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_775_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_775_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_776_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_776_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_777_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_777_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_778_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_778_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_779_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_779_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_780_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_780_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_781_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_781_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_782_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_782_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_783_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_783_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_784_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_784_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_785_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_785_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_786_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_786_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_787_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_787_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_788_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_788_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_789_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_789_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_790_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_790_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_791_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_791_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_792_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_792_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_793_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_793_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_794_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_794_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_795_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_795_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_796_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_796_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_797_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_797_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_798_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_798_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_799_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_799_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_800_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_800_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_801_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_801_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_802_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_802_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_803_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_803_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_804_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_804_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_805_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_805_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_806_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_806_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_807_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_807_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_808_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_808_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_809_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_809_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_810_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_810_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_811_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_811_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_812_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_812_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_813_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_813_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_814_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_814_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_815_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_815_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_816_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_816_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_817_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_817_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_818_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_818_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_819_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_819_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_820_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_820_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_821_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_821_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_822_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_822_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_823_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_823_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_824_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_824_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_825_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_825_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_826_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_826_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_827_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_827_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_828_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_828_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_829_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_829_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_830_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_830_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_831_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_831_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_832_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_832_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_833_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_833_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_834_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_834_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_835_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_835_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_836_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_836_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_837_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_837_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_838_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_838_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_839_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_839_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_840_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_840_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_841_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_841_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_842_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_842_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_843_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_843_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_844_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_844_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_845_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_845_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_846_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_846_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_847_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_847_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_848_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_848_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_849_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_849_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_850_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_850_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_851_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_851_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_852_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_852_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_853_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_853_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_854_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_854_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_855_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_855_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_856_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_856_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_857_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_857_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_858_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_858_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_859_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_859_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_860_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_860_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_861_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_861_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_862_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_862_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_863_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_863_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_864_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_864_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_865_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_865_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_866_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_866_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_867_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_867_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_868_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_868_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_869_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_869_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_870_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_870_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_871_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_871_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_872_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_872_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_873_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_873_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_874_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_874_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_875_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_875_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_876_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_876_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_877_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_877_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_878_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_878_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_879_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_879_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_880_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_880_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_881_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_881_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_882_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_882_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_883_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_883_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_884_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_884_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_885_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_885_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_886_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_886_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_887_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_887_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_888_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_888_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_889_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_889_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_890_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_890_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_891_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_891_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_892_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_892_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_893_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_893_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_894_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_894_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_895_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_895_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_896_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_896_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_897_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_897_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_898_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_898_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_899_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_899_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_900_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_900_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_901_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_901_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_902_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_902_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_903_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_903_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_904_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_904_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_905_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_905_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_906_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_906_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_907_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_907_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_908_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_908_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_909_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_909_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_910_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_910_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_911_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_911_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_912_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_912_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_913_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_913_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_914_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_914_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_915_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_915_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_916_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_916_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_917_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_917_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_918_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_918_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_919_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_919_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_920_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_920_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_921_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_921_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_922_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_922_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_923_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_923_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_924_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_924_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_925_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_925_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_926_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_926_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_927_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_927_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_928_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_928_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_929_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_929_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_930_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_930_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_931_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_931_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_932_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_932_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_933_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_933_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_934_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_934_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_935_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_935_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_936_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_936_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_937_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_937_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_938_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_938_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_939_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_939_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_940_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_940_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_941_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_941_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_942_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_942_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_943_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_943_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_944_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_944_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_945_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_945_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_946_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_946_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_947_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_947_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_948_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_948_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_949_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_949_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_950_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_950_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_951_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_951_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_952_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_952_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_953_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_953_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_954_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_954_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_955_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_955_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_956_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_956_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_957_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_957_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_958_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_958_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_959_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_959_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_960_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_960_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_961_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_961_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_962_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_962_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_963_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_963_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_964_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_964_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_965_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_965_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_966_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_966_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_967_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_967_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_968_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_968_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_969_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_969_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_970_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_970_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_971_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_971_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_972_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_972_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_973_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_973_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_974_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_974_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_975_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_975_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_976_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_976_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_977_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_977_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_978_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_978_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_979_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_979_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_980_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_980_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_981_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_981_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_982_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_982_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_983_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_983_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_984_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_984_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_985_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_985_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_986_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_986_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_987_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_987_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_988_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_988_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_989_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_989_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_990_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_990_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_991_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_991_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_992_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_992_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_993_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_993_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_994_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_994_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_995_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_995_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_996_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_996_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_997_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_997_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_998_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_998_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_999_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_999_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1000_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1000_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1001_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1001_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1002_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1002_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1003_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1003_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1004_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1004_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1005_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1005_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1006_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1006_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1007_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1007_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1008_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1008_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1009_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1009_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1010_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1010_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1011_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1011_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1012_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1012_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1013_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1013_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1014_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1014_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1015_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1015_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1016_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1016_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1017_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1017_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1018_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1018_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1019_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1019_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1020_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1020_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1021_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1021_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1022_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1022_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1023_0; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  reg  r_1023_1; // @[src/main/scala/gemmini/Mesh.scala 112:41]
  Tile mesh_0_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_0_clock),
    .io_in_a_0(mesh_0_0_io_in_a_0),
    .io_in_a_1(mesh_0_0_io_in_a_1),
    .io_in_b_0(mesh_0_0_io_in_b_0),
    .io_in_b_1(mesh_0_0_io_in_b_1),
    .io_in_d_0(mesh_0_0_io_in_d_0),
    .io_in_d_1(mesh_0_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_0_io_in_control_1_shift),
    .io_in_id_0(mesh_0_0_io_in_id_0),
    .io_in_id_1(mesh_0_0_io_in_id_1),
    .io_in_last_0(mesh_0_0_io_in_last_0),
    .io_in_last_1(mesh_0_0_io_in_last_1),
    .io_out_a_0(mesh_0_0_io_out_a_0),
    .io_out_a_1(mesh_0_0_io_out_a_1),
    .io_out_c_0(mesh_0_0_io_out_c_0),
    .io_out_c_1(mesh_0_0_io_out_c_1),
    .io_out_b_0(mesh_0_0_io_out_b_0),
    .io_out_b_1(mesh_0_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_0_io_out_control_1_shift),
    .io_out_id_0(mesh_0_0_io_out_id_0),
    .io_out_id_1(mesh_0_0_io_out_id_1),
    .io_out_last_0(mesh_0_0_io_out_last_0),
    .io_out_last_1(mesh_0_0_io_out_last_1),
    .io_in_valid_0(mesh_0_0_io_in_valid_0),
    .io_in_valid_1(mesh_0_0_io_in_valid_1),
    .io_out_valid_0(mesh_0_0_io_out_valid_0),
    .io_out_valid_1(mesh_0_0_io_out_valid_1)
  );
  Tile mesh_0_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_1_clock),
    .io_in_a_0(mesh_0_1_io_in_a_0),
    .io_in_a_1(mesh_0_1_io_in_a_1),
    .io_in_b_0(mesh_0_1_io_in_b_0),
    .io_in_b_1(mesh_0_1_io_in_b_1),
    .io_in_d_0(mesh_0_1_io_in_d_0),
    .io_in_d_1(mesh_0_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_1_io_in_control_1_shift),
    .io_in_id_0(mesh_0_1_io_in_id_0),
    .io_in_id_1(mesh_0_1_io_in_id_1),
    .io_in_last_0(mesh_0_1_io_in_last_0),
    .io_in_last_1(mesh_0_1_io_in_last_1),
    .io_out_a_0(mesh_0_1_io_out_a_0),
    .io_out_a_1(mesh_0_1_io_out_a_1),
    .io_out_c_0(mesh_0_1_io_out_c_0),
    .io_out_c_1(mesh_0_1_io_out_c_1),
    .io_out_b_0(mesh_0_1_io_out_b_0),
    .io_out_b_1(mesh_0_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_1_io_out_control_1_shift),
    .io_out_id_0(mesh_0_1_io_out_id_0),
    .io_out_id_1(mesh_0_1_io_out_id_1),
    .io_out_last_0(mesh_0_1_io_out_last_0),
    .io_out_last_1(mesh_0_1_io_out_last_1),
    .io_in_valid_0(mesh_0_1_io_in_valid_0),
    .io_in_valid_1(mesh_0_1_io_in_valid_1),
    .io_out_valid_0(mesh_0_1_io_out_valid_0),
    .io_out_valid_1(mesh_0_1_io_out_valid_1)
  );
  Tile mesh_0_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_2_clock),
    .io_in_a_0(mesh_0_2_io_in_a_0),
    .io_in_a_1(mesh_0_2_io_in_a_1),
    .io_in_b_0(mesh_0_2_io_in_b_0),
    .io_in_b_1(mesh_0_2_io_in_b_1),
    .io_in_d_0(mesh_0_2_io_in_d_0),
    .io_in_d_1(mesh_0_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_2_io_in_control_1_shift),
    .io_in_id_0(mesh_0_2_io_in_id_0),
    .io_in_id_1(mesh_0_2_io_in_id_1),
    .io_in_last_0(mesh_0_2_io_in_last_0),
    .io_in_last_1(mesh_0_2_io_in_last_1),
    .io_out_a_0(mesh_0_2_io_out_a_0),
    .io_out_a_1(mesh_0_2_io_out_a_1),
    .io_out_c_0(mesh_0_2_io_out_c_0),
    .io_out_c_1(mesh_0_2_io_out_c_1),
    .io_out_b_0(mesh_0_2_io_out_b_0),
    .io_out_b_1(mesh_0_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_2_io_out_control_1_shift),
    .io_out_id_0(mesh_0_2_io_out_id_0),
    .io_out_id_1(mesh_0_2_io_out_id_1),
    .io_out_last_0(mesh_0_2_io_out_last_0),
    .io_out_last_1(mesh_0_2_io_out_last_1),
    .io_in_valid_0(mesh_0_2_io_in_valid_0),
    .io_in_valid_1(mesh_0_2_io_in_valid_1),
    .io_out_valid_0(mesh_0_2_io_out_valid_0),
    .io_out_valid_1(mesh_0_2_io_out_valid_1)
  );
  Tile mesh_0_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_3_clock),
    .io_in_a_0(mesh_0_3_io_in_a_0),
    .io_in_a_1(mesh_0_3_io_in_a_1),
    .io_in_b_0(mesh_0_3_io_in_b_0),
    .io_in_b_1(mesh_0_3_io_in_b_1),
    .io_in_d_0(mesh_0_3_io_in_d_0),
    .io_in_d_1(mesh_0_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_3_io_in_control_1_shift),
    .io_in_id_0(mesh_0_3_io_in_id_0),
    .io_in_id_1(mesh_0_3_io_in_id_1),
    .io_in_last_0(mesh_0_3_io_in_last_0),
    .io_in_last_1(mesh_0_3_io_in_last_1),
    .io_out_a_0(mesh_0_3_io_out_a_0),
    .io_out_a_1(mesh_0_3_io_out_a_1),
    .io_out_c_0(mesh_0_3_io_out_c_0),
    .io_out_c_1(mesh_0_3_io_out_c_1),
    .io_out_b_0(mesh_0_3_io_out_b_0),
    .io_out_b_1(mesh_0_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_3_io_out_control_1_shift),
    .io_out_id_0(mesh_0_3_io_out_id_0),
    .io_out_id_1(mesh_0_3_io_out_id_1),
    .io_out_last_0(mesh_0_3_io_out_last_0),
    .io_out_last_1(mesh_0_3_io_out_last_1),
    .io_in_valid_0(mesh_0_3_io_in_valid_0),
    .io_in_valid_1(mesh_0_3_io_in_valid_1),
    .io_out_valid_0(mesh_0_3_io_out_valid_0),
    .io_out_valid_1(mesh_0_3_io_out_valid_1)
  );
  Tile mesh_0_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_4_clock),
    .io_in_a_0(mesh_0_4_io_in_a_0),
    .io_in_a_1(mesh_0_4_io_in_a_1),
    .io_in_b_0(mesh_0_4_io_in_b_0),
    .io_in_b_1(mesh_0_4_io_in_b_1),
    .io_in_d_0(mesh_0_4_io_in_d_0),
    .io_in_d_1(mesh_0_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_4_io_in_control_1_shift),
    .io_in_id_0(mesh_0_4_io_in_id_0),
    .io_in_id_1(mesh_0_4_io_in_id_1),
    .io_in_last_0(mesh_0_4_io_in_last_0),
    .io_in_last_1(mesh_0_4_io_in_last_1),
    .io_out_a_0(mesh_0_4_io_out_a_0),
    .io_out_a_1(mesh_0_4_io_out_a_1),
    .io_out_c_0(mesh_0_4_io_out_c_0),
    .io_out_c_1(mesh_0_4_io_out_c_1),
    .io_out_b_0(mesh_0_4_io_out_b_0),
    .io_out_b_1(mesh_0_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_4_io_out_control_1_shift),
    .io_out_id_0(mesh_0_4_io_out_id_0),
    .io_out_id_1(mesh_0_4_io_out_id_1),
    .io_out_last_0(mesh_0_4_io_out_last_0),
    .io_out_last_1(mesh_0_4_io_out_last_1),
    .io_in_valid_0(mesh_0_4_io_in_valid_0),
    .io_in_valid_1(mesh_0_4_io_in_valid_1),
    .io_out_valid_0(mesh_0_4_io_out_valid_0),
    .io_out_valid_1(mesh_0_4_io_out_valid_1)
  );
  Tile mesh_0_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_5_clock),
    .io_in_a_0(mesh_0_5_io_in_a_0),
    .io_in_a_1(mesh_0_5_io_in_a_1),
    .io_in_b_0(mesh_0_5_io_in_b_0),
    .io_in_b_1(mesh_0_5_io_in_b_1),
    .io_in_d_0(mesh_0_5_io_in_d_0),
    .io_in_d_1(mesh_0_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_5_io_in_control_1_shift),
    .io_in_id_0(mesh_0_5_io_in_id_0),
    .io_in_id_1(mesh_0_5_io_in_id_1),
    .io_in_last_0(mesh_0_5_io_in_last_0),
    .io_in_last_1(mesh_0_5_io_in_last_1),
    .io_out_a_0(mesh_0_5_io_out_a_0),
    .io_out_a_1(mesh_0_5_io_out_a_1),
    .io_out_c_0(mesh_0_5_io_out_c_0),
    .io_out_c_1(mesh_0_5_io_out_c_1),
    .io_out_b_0(mesh_0_5_io_out_b_0),
    .io_out_b_1(mesh_0_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_5_io_out_control_1_shift),
    .io_out_id_0(mesh_0_5_io_out_id_0),
    .io_out_id_1(mesh_0_5_io_out_id_1),
    .io_out_last_0(mesh_0_5_io_out_last_0),
    .io_out_last_1(mesh_0_5_io_out_last_1),
    .io_in_valid_0(mesh_0_5_io_in_valid_0),
    .io_in_valid_1(mesh_0_5_io_in_valid_1),
    .io_out_valid_0(mesh_0_5_io_out_valid_0),
    .io_out_valid_1(mesh_0_5_io_out_valid_1)
  );
  Tile mesh_0_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_6_clock),
    .io_in_a_0(mesh_0_6_io_in_a_0),
    .io_in_a_1(mesh_0_6_io_in_a_1),
    .io_in_b_0(mesh_0_6_io_in_b_0),
    .io_in_b_1(mesh_0_6_io_in_b_1),
    .io_in_d_0(mesh_0_6_io_in_d_0),
    .io_in_d_1(mesh_0_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_6_io_in_control_1_shift),
    .io_in_id_0(mesh_0_6_io_in_id_0),
    .io_in_id_1(mesh_0_6_io_in_id_1),
    .io_in_last_0(mesh_0_6_io_in_last_0),
    .io_in_last_1(mesh_0_6_io_in_last_1),
    .io_out_a_0(mesh_0_6_io_out_a_0),
    .io_out_a_1(mesh_0_6_io_out_a_1),
    .io_out_c_0(mesh_0_6_io_out_c_0),
    .io_out_c_1(mesh_0_6_io_out_c_1),
    .io_out_b_0(mesh_0_6_io_out_b_0),
    .io_out_b_1(mesh_0_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_6_io_out_control_1_shift),
    .io_out_id_0(mesh_0_6_io_out_id_0),
    .io_out_id_1(mesh_0_6_io_out_id_1),
    .io_out_last_0(mesh_0_6_io_out_last_0),
    .io_out_last_1(mesh_0_6_io_out_last_1),
    .io_in_valid_0(mesh_0_6_io_in_valid_0),
    .io_in_valid_1(mesh_0_6_io_in_valid_1),
    .io_out_valid_0(mesh_0_6_io_out_valid_0),
    .io_out_valid_1(mesh_0_6_io_out_valid_1)
  );
  Tile mesh_0_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_7_clock),
    .io_in_a_0(mesh_0_7_io_in_a_0),
    .io_in_a_1(mesh_0_7_io_in_a_1),
    .io_in_b_0(mesh_0_7_io_in_b_0),
    .io_in_b_1(mesh_0_7_io_in_b_1),
    .io_in_d_0(mesh_0_7_io_in_d_0),
    .io_in_d_1(mesh_0_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_7_io_in_control_1_shift),
    .io_in_id_0(mesh_0_7_io_in_id_0),
    .io_in_id_1(mesh_0_7_io_in_id_1),
    .io_in_last_0(mesh_0_7_io_in_last_0),
    .io_in_last_1(mesh_0_7_io_in_last_1),
    .io_out_a_0(mesh_0_7_io_out_a_0),
    .io_out_a_1(mesh_0_7_io_out_a_1),
    .io_out_c_0(mesh_0_7_io_out_c_0),
    .io_out_c_1(mesh_0_7_io_out_c_1),
    .io_out_b_0(mesh_0_7_io_out_b_0),
    .io_out_b_1(mesh_0_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_7_io_out_control_1_shift),
    .io_out_id_0(mesh_0_7_io_out_id_0),
    .io_out_id_1(mesh_0_7_io_out_id_1),
    .io_out_last_0(mesh_0_7_io_out_last_0),
    .io_out_last_1(mesh_0_7_io_out_last_1),
    .io_in_valid_0(mesh_0_7_io_in_valid_0),
    .io_in_valid_1(mesh_0_7_io_in_valid_1),
    .io_out_valid_0(mesh_0_7_io_out_valid_0),
    .io_out_valid_1(mesh_0_7_io_out_valid_1)
  );
  Tile mesh_0_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_8_clock),
    .io_in_a_0(mesh_0_8_io_in_a_0),
    .io_in_a_1(mesh_0_8_io_in_a_1),
    .io_in_b_0(mesh_0_8_io_in_b_0),
    .io_in_b_1(mesh_0_8_io_in_b_1),
    .io_in_d_0(mesh_0_8_io_in_d_0),
    .io_in_d_1(mesh_0_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_8_io_in_control_1_shift),
    .io_in_id_0(mesh_0_8_io_in_id_0),
    .io_in_id_1(mesh_0_8_io_in_id_1),
    .io_in_last_0(mesh_0_8_io_in_last_0),
    .io_in_last_1(mesh_0_8_io_in_last_1),
    .io_out_a_0(mesh_0_8_io_out_a_0),
    .io_out_a_1(mesh_0_8_io_out_a_1),
    .io_out_c_0(mesh_0_8_io_out_c_0),
    .io_out_c_1(mesh_0_8_io_out_c_1),
    .io_out_b_0(mesh_0_8_io_out_b_0),
    .io_out_b_1(mesh_0_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_8_io_out_control_1_shift),
    .io_out_id_0(mesh_0_8_io_out_id_0),
    .io_out_id_1(mesh_0_8_io_out_id_1),
    .io_out_last_0(mesh_0_8_io_out_last_0),
    .io_out_last_1(mesh_0_8_io_out_last_1),
    .io_in_valid_0(mesh_0_8_io_in_valid_0),
    .io_in_valid_1(mesh_0_8_io_in_valid_1),
    .io_out_valid_0(mesh_0_8_io_out_valid_0),
    .io_out_valid_1(mesh_0_8_io_out_valid_1)
  );
  Tile mesh_0_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_9_clock),
    .io_in_a_0(mesh_0_9_io_in_a_0),
    .io_in_a_1(mesh_0_9_io_in_a_1),
    .io_in_b_0(mesh_0_9_io_in_b_0),
    .io_in_b_1(mesh_0_9_io_in_b_1),
    .io_in_d_0(mesh_0_9_io_in_d_0),
    .io_in_d_1(mesh_0_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_9_io_in_control_1_shift),
    .io_in_id_0(mesh_0_9_io_in_id_0),
    .io_in_id_1(mesh_0_9_io_in_id_1),
    .io_in_last_0(mesh_0_9_io_in_last_0),
    .io_in_last_1(mesh_0_9_io_in_last_1),
    .io_out_a_0(mesh_0_9_io_out_a_0),
    .io_out_a_1(mesh_0_9_io_out_a_1),
    .io_out_c_0(mesh_0_9_io_out_c_0),
    .io_out_c_1(mesh_0_9_io_out_c_1),
    .io_out_b_0(mesh_0_9_io_out_b_0),
    .io_out_b_1(mesh_0_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_9_io_out_control_1_shift),
    .io_out_id_0(mesh_0_9_io_out_id_0),
    .io_out_id_1(mesh_0_9_io_out_id_1),
    .io_out_last_0(mesh_0_9_io_out_last_0),
    .io_out_last_1(mesh_0_9_io_out_last_1),
    .io_in_valid_0(mesh_0_9_io_in_valid_0),
    .io_in_valid_1(mesh_0_9_io_in_valid_1),
    .io_out_valid_0(mesh_0_9_io_out_valid_0),
    .io_out_valid_1(mesh_0_9_io_out_valid_1)
  );
  Tile mesh_0_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_10_clock),
    .io_in_a_0(mesh_0_10_io_in_a_0),
    .io_in_a_1(mesh_0_10_io_in_a_1),
    .io_in_b_0(mesh_0_10_io_in_b_0),
    .io_in_b_1(mesh_0_10_io_in_b_1),
    .io_in_d_0(mesh_0_10_io_in_d_0),
    .io_in_d_1(mesh_0_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_10_io_in_control_1_shift),
    .io_in_id_0(mesh_0_10_io_in_id_0),
    .io_in_id_1(mesh_0_10_io_in_id_1),
    .io_in_last_0(mesh_0_10_io_in_last_0),
    .io_in_last_1(mesh_0_10_io_in_last_1),
    .io_out_a_0(mesh_0_10_io_out_a_0),
    .io_out_a_1(mesh_0_10_io_out_a_1),
    .io_out_c_0(mesh_0_10_io_out_c_0),
    .io_out_c_1(mesh_0_10_io_out_c_1),
    .io_out_b_0(mesh_0_10_io_out_b_0),
    .io_out_b_1(mesh_0_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_10_io_out_control_1_shift),
    .io_out_id_0(mesh_0_10_io_out_id_0),
    .io_out_id_1(mesh_0_10_io_out_id_1),
    .io_out_last_0(mesh_0_10_io_out_last_0),
    .io_out_last_1(mesh_0_10_io_out_last_1),
    .io_in_valid_0(mesh_0_10_io_in_valid_0),
    .io_in_valid_1(mesh_0_10_io_in_valid_1),
    .io_out_valid_0(mesh_0_10_io_out_valid_0),
    .io_out_valid_1(mesh_0_10_io_out_valid_1)
  );
  Tile mesh_0_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_11_clock),
    .io_in_a_0(mesh_0_11_io_in_a_0),
    .io_in_a_1(mesh_0_11_io_in_a_1),
    .io_in_b_0(mesh_0_11_io_in_b_0),
    .io_in_b_1(mesh_0_11_io_in_b_1),
    .io_in_d_0(mesh_0_11_io_in_d_0),
    .io_in_d_1(mesh_0_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_11_io_in_control_1_shift),
    .io_in_id_0(mesh_0_11_io_in_id_0),
    .io_in_id_1(mesh_0_11_io_in_id_1),
    .io_in_last_0(mesh_0_11_io_in_last_0),
    .io_in_last_1(mesh_0_11_io_in_last_1),
    .io_out_a_0(mesh_0_11_io_out_a_0),
    .io_out_a_1(mesh_0_11_io_out_a_1),
    .io_out_c_0(mesh_0_11_io_out_c_0),
    .io_out_c_1(mesh_0_11_io_out_c_1),
    .io_out_b_0(mesh_0_11_io_out_b_0),
    .io_out_b_1(mesh_0_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_11_io_out_control_1_shift),
    .io_out_id_0(mesh_0_11_io_out_id_0),
    .io_out_id_1(mesh_0_11_io_out_id_1),
    .io_out_last_0(mesh_0_11_io_out_last_0),
    .io_out_last_1(mesh_0_11_io_out_last_1),
    .io_in_valid_0(mesh_0_11_io_in_valid_0),
    .io_in_valid_1(mesh_0_11_io_in_valid_1),
    .io_out_valid_0(mesh_0_11_io_out_valid_0),
    .io_out_valid_1(mesh_0_11_io_out_valid_1)
  );
  Tile mesh_0_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_12_clock),
    .io_in_a_0(mesh_0_12_io_in_a_0),
    .io_in_a_1(mesh_0_12_io_in_a_1),
    .io_in_b_0(mesh_0_12_io_in_b_0),
    .io_in_b_1(mesh_0_12_io_in_b_1),
    .io_in_d_0(mesh_0_12_io_in_d_0),
    .io_in_d_1(mesh_0_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_12_io_in_control_1_shift),
    .io_in_id_0(mesh_0_12_io_in_id_0),
    .io_in_id_1(mesh_0_12_io_in_id_1),
    .io_in_last_0(mesh_0_12_io_in_last_0),
    .io_in_last_1(mesh_0_12_io_in_last_1),
    .io_out_a_0(mesh_0_12_io_out_a_0),
    .io_out_a_1(mesh_0_12_io_out_a_1),
    .io_out_c_0(mesh_0_12_io_out_c_0),
    .io_out_c_1(mesh_0_12_io_out_c_1),
    .io_out_b_0(mesh_0_12_io_out_b_0),
    .io_out_b_1(mesh_0_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_12_io_out_control_1_shift),
    .io_out_id_0(mesh_0_12_io_out_id_0),
    .io_out_id_1(mesh_0_12_io_out_id_1),
    .io_out_last_0(mesh_0_12_io_out_last_0),
    .io_out_last_1(mesh_0_12_io_out_last_1),
    .io_in_valid_0(mesh_0_12_io_in_valid_0),
    .io_in_valid_1(mesh_0_12_io_in_valid_1),
    .io_out_valid_0(mesh_0_12_io_out_valid_0),
    .io_out_valid_1(mesh_0_12_io_out_valid_1)
  );
  Tile mesh_0_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_13_clock),
    .io_in_a_0(mesh_0_13_io_in_a_0),
    .io_in_a_1(mesh_0_13_io_in_a_1),
    .io_in_b_0(mesh_0_13_io_in_b_0),
    .io_in_b_1(mesh_0_13_io_in_b_1),
    .io_in_d_0(mesh_0_13_io_in_d_0),
    .io_in_d_1(mesh_0_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_13_io_in_control_1_shift),
    .io_in_id_0(mesh_0_13_io_in_id_0),
    .io_in_id_1(mesh_0_13_io_in_id_1),
    .io_in_last_0(mesh_0_13_io_in_last_0),
    .io_in_last_1(mesh_0_13_io_in_last_1),
    .io_out_a_0(mesh_0_13_io_out_a_0),
    .io_out_a_1(mesh_0_13_io_out_a_1),
    .io_out_c_0(mesh_0_13_io_out_c_0),
    .io_out_c_1(mesh_0_13_io_out_c_1),
    .io_out_b_0(mesh_0_13_io_out_b_0),
    .io_out_b_1(mesh_0_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_13_io_out_control_1_shift),
    .io_out_id_0(mesh_0_13_io_out_id_0),
    .io_out_id_1(mesh_0_13_io_out_id_1),
    .io_out_last_0(mesh_0_13_io_out_last_0),
    .io_out_last_1(mesh_0_13_io_out_last_1),
    .io_in_valid_0(mesh_0_13_io_in_valid_0),
    .io_in_valid_1(mesh_0_13_io_in_valid_1),
    .io_out_valid_0(mesh_0_13_io_out_valid_0),
    .io_out_valid_1(mesh_0_13_io_out_valid_1)
  );
  Tile mesh_0_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_14_clock),
    .io_in_a_0(mesh_0_14_io_in_a_0),
    .io_in_a_1(mesh_0_14_io_in_a_1),
    .io_in_b_0(mesh_0_14_io_in_b_0),
    .io_in_b_1(mesh_0_14_io_in_b_1),
    .io_in_d_0(mesh_0_14_io_in_d_0),
    .io_in_d_1(mesh_0_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_14_io_in_control_1_shift),
    .io_in_id_0(mesh_0_14_io_in_id_0),
    .io_in_id_1(mesh_0_14_io_in_id_1),
    .io_in_last_0(mesh_0_14_io_in_last_0),
    .io_in_last_1(mesh_0_14_io_in_last_1),
    .io_out_a_0(mesh_0_14_io_out_a_0),
    .io_out_a_1(mesh_0_14_io_out_a_1),
    .io_out_c_0(mesh_0_14_io_out_c_0),
    .io_out_c_1(mesh_0_14_io_out_c_1),
    .io_out_b_0(mesh_0_14_io_out_b_0),
    .io_out_b_1(mesh_0_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_14_io_out_control_1_shift),
    .io_out_id_0(mesh_0_14_io_out_id_0),
    .io_out_id_1(mesh_0_14_io_out_id_1),
    .io_out_last_0(mesh_0_14_io_out_last_0),
    .io_out_last_1(mesh_0_14_io_out_last_1),
    .io_in_valid_0(mesh_0_14_io_in_valid_0),
    .io_in_valid_1(mesh_0_14_io_in_valid_1),
    .io_out_valid_0(mesh_0_14_io_out_valid_0),
    .io_out_valid_1(mesh_0_14_io_out_valid_1)
  );
  Tile mesh_0_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_0_15_clock),
    .io_in_a_0(mesh_0_15_io_in_a_0),
    .io_in_a_1(mesh_0_15_io_in_a_1),
    .io_in_b_0(mesh_0_15_io_in_b_0),
    .io_in_b_1(mesh_0_15_io_in_b_1),
    .io_in_d_0(mesh_0_15_io_in_d_0),
    .io_in_d_1(mesh_0_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_15_io_in_control_1_shift),
    .io_in_id_0(mesh_0_15_io_in_id_0),
    .io_in_id_1(mesh_0_15_io_in_id_1),
    .io_in_last_0(mesh_0_15_io_in_last_0),
    .io_in_last_1(mesh_0_15_io_in_last_1),
    .io_out_a_0(mesh_0_15_io_out_a_0),
    .io_out_a_1(mesh_0_15_io_out_a_1),
    .io_out_c_0(mesh_0_15_io_out_c_0),
    .io_out_c_1(mesh_0_15_io_out_c_1),
    .io_out_b_0(mesh_0_15_io_out_b_0),
    .io_out_b_1(mesh_0_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_15_io_out_control_1_shift),
    .io_out_id_0(mesh_0_15_io_out_id_0),
    .io_out_id_1(mesh_0_15_io_out_id_1),
    .io_out_last_0(mesh_0_15_io_out_last_0),
    .io_out_last_1(mesh_0_15_io_out_last_1),
    .io_in_valid_0(mesh_0_15_io_in_valid_0),
    .io_in_valid_1(mesh_0_15_io_in_valid_1),
    .io_out_valid_0(mesh_0_15_io_out_valid_0),
    .io_out_valid_1(mesh_0_15_io_out_valid_1)
  );
  Tile mesh_1_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_0_clock),
    .io_in_a_0(mesh_1_0_io_in_a_0),
    .io_in_a_1(mesh_1_0_io_in_a_1),
    .io_in_b_0(mesh_1_0_io_in_b_0),
    .io_in_b_1(mesh_1_0_io_in_b_1),
    .io_in_d_0(mesh_1_0_io_in_d_0),
    .io_in_d_1(mesh_1_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_0_io_in_control_1_shift),
    .io_in_id_0(mesh_1_0_io_in_id_0),
    .io_in_id_1(mesh_1_0_io_in_id_1),
    .io_in_last_0(mesh_1_0_io_in_last_0),
    .io_in_last_1(mesh_1_0_io_in_last_1),
    .io_out_a_0(mesh_1_0_io_out_a_0),
    .io_out_a_1(mesh_1_0_io_out_a_1),
    .io_out_c_0(mesh_1_0_io_out_c_0),
    .io_out_c_1(mesh_1_0_io_out_c_1),
    .io_out_b_0(mesh_1_0_io_out_b_0),
    .io_out_b_1(mesh_1_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_0_io_out_control_1_shift),
    .io_out_id_0(mesh_1_0_io_out_id_0),
    .io_out_id_1(mesh_1_0_io_out_id_1),
    .io_out_last_0(mesh_1_0_io_out_last_0),
    .io_out_last_1(mesh_1_0_io_out_last_1),
    .io_in_valid_0(mesh_1_0_io_in_valid_0),
    .io_in_valid_1(mesh_1_0_io_in_valid_1),
    .io_out_valid_0(mesh_1_0_io_out_valid_0),
    .io_out_valid_1(mesh_1_0_io_out_valid_1)
  );
  Tile mesh_1_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_1_clock),
    .io_in_a_0(mesh_1_1_io_in_a_0),
    .io_in_a_1(mesh_1_1_io_in_a_1),
    .io_in_b_0(mesh_1_1_io_in_b_0),
    .io_in_b_1(mesh_1_1_io_in_b_1),
    .io_in_d_0(mesh_1_1_io_in_d_0),
    .io_in_d_1(mesh_1_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_1_io_in_control_1_shift),
    .io_in_id_0(mesh_1_1_io_in_id_0),
    .io_in_id_1(mesh_1_1_io_in_id_1),
    .io_in_last_0(mesh_1_1_io_in_last_0),
    .io_in_last_1(mesh_1_1_io_in_last_1),
    .io_out_a_0(mesh_1_1_io_out_a_0),
    .io_out_a_1(mesh_1_1_io_out_a_1),
    .io_out_c_0(mesh_1_1_io_out_c_0),
    .io_out_c_1(mesh_1_1_io_out_c_1),
    .io_out_b_0(mesh_1_1_io_out_b_0),
    .io_out_b_1(mesh_1_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_1_io_out_control_1_shift),
    .io_out_id_0(mesh_1_1_io_out_id_0),
    .io_out_id_1(mesh_1_1_io_out_id_1),
    .io_out_last_0(mesh_1_1_io_out_last_0),
    .io_out_last_1(mesh_1_1_io_out_last_1),
    .io_in_valid_0(mesh_1_1_io_in_valid_0),
    .io_in_valid_1(mesh_1_1_io_in_valid_1),
    .io_out_valid_0(mesh_1_1_io_out_valid_0),
    .io_out_valid_1(mesh_1_1_io_out_valid_1)
  );
  Tile mesh_1_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_2_clock),
    .io_in_a_0(mesh_1_2_io_in_a_0),
    .io_in_a_1(mesh_1_2_io_in_a_1),
    .io_in_b_0(mesh_1_2_io_in_b_0),
    .io_in_b_1(mesh_1_2_io_in_b_1),
    .io_in_d_0(mesh_1_2_io_in_d_0),
    .io_in_d_1(mesh_1_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_2_io_in_control_1_shift),
    .io_in_id_0(mesh_1_2_io_in_id_0),
    .io_in_id_1(mesh_1_2_io_in_id_1),
    .io_in_last_0(mesh_1_2_io_in_last_0),
    .io_in_last_1(mesh_1_2_io_in_last_1),
    .io_out_a_0(mesh_1_2_io_out_a_0),
    .io_out_a_1(mesh_1_2_io_out_a_1),
    .io_out_c_0(mesh_1_2_io_out_c_0),
    .io_out_c_1(mesh_1_2_io_out_c_1),
    .io_out_b_0(mesh_1_2_io_out_b_0),
    .io_out_b_1(mesh_1_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_2_io_out_control_1_shift),
    .io_out_id_0(mesh_1_2_io_out_id_0),
    .io_out_id_1(mesh_1_2_io_out_id_1),
    .io_out_last_0(mesh_1_2_io_out_last_0),
    .io_out_last_1(mesh_1_2_io_out_last_1),
    .io_in_valid_0(mesh_1_2_io_in_valid_0),
    .io_in_valid_1(mesh_1_2_io_in_valid_1),
    .io_out_valid_0(mesh_1_2_io_out_valid_0),
    .io_out_valid_1(mesh_1_2_io_out_valid_1)
  );
  Tile mesh_1_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_3_clock),
    .io_in_a_0(mesh_1_3_io_in_a_0),
    .io_in_a_1(mesh_1_3_io_in_a_1),
    .io_in_b_0(mesh_1_3_io_in_b_0),
    .io_in_b_1(mesh_1_3_io_in_b_1),
    .io_in_d_0(mesh_1_3_io_in_d_0),
    .io_in_d_1(mesh_1_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_3_io_in_control_1_shift),
    .io_in_id_0(mesh_1_3_io_in_id_0),
    .io_in_id_1(mesh_1_3_io_in_id_1),
    .io_in_last_0(mesh_1_3_io_in_last_0),
    .io_in_last_1(mesh_1_3_io_in_last_1),
    .io_out_a_0(mesh_1_3_io_out_a_0),
    .io_out_a_1(mesh_1_3_io_out_a_1),
    .io_out_c_0(mesh_1_3_io_out_c_0),
    .io_out_c_1(mesh_1_3_io_out_c_1),
    .io_out_b_0(mesh_1_3_io_out_b_0),
    .io_out_b_1(mesh_1_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_3_io_out_control_1_shift),
    .io_out_id_0(mesh_1_3_io_out_id_0),
    .io_out_id_1(mesh_1_3_io_out_id_1),
    .io_out_last_0(mesh_1_3_io_out_last_0),
    .io_out_last_1(mesh_1_3_io_out_last_1),
    .io_in_valid_0(mesh_1_3_io_in_valid_0),
    .io_in_valid_1(mesh_1_3_io_in_valid_1),
    .io_out_valid_0(mesh_1_3_io_out_valid_0),
    .io_out_valid_1(mesh_1_3_io_out_valid_1)
  );
  Tile mesh_1_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_4_clock),
    .io_in_a_0(mesh_1_4_io_in_a_0),
    .io_in_a_1(mesh_1_4_io_in_a_1),
    .io_in_b_0(mesh_1_4_io_in_b_0),
    .io_in_b_1(mesh_1_4_io_in_b_1),
    .io_in_d_0(mesh_1_4_io_in_d_0),
    .io_in_d_1(mesh_1_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_4_io_in_control_1_shift),
    .io_in_id_0(mesh_1_4_io_in_id_0),
    .io_in_id_1(mesh_1_4_io_in_id_1),
    .io_in_last_0(mesh_1_4_io_in_last_0),
    .io_in_last_1(mesh_1_4_io_in_last_1),
    .io_out_a_0(mesh_1_4_io_out_a_0),
    .io_out_a_1(mesh_1_4_io_out_a_1),
    .io_out_c_0(mesh_1_4_io_out_c_0),
    .io_out_c_1(mesh_1_4_io_out_c_1),
    .io_out_b_0(mesh_1_4_io_out_b_0),
    .io_out_b_1(mesh_1_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_4_io_out_control_1_shift),
    .io_out_id_0(mesh_1_4_io_out_id_0),
    .io_out_id_1(mesh_1_4_io_out_id_1),
    .io_out_last_0(mesh_1_4_io_out_last_0),
    .io_out_last_1(mesh_1_4_io_out_last_1),
    .io_in_valid_0(mesh_1_4_io_in_valid_0),
    .io_in_valid_1(mesh_1_4_io_in_valid_1),
    .io_out_valid_0(mesh_1_4_io_out_valid_0),
    .io_out_valid_1(mesh_1_4_io_out_valid_1)
  );
  Tile mesh_1_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_5_clock),
    .io_in_a_0(mesh_1_5_io_in_a_0),
    .io_in_a_1(mesh_1_5_io_in_a_1),
    .io_in_b_0(mesh_1_5_io_in_b_0),
    .io_in_b_1(mesh_1_5_io_in_b_1),
    .io_in_d_0(mesh_1_5_io_in_d_0),
    .io_in_d_1(mesh_1_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_5_io_in_control_1_shift),
    .io_in_id_0(mesh_1_5_io_in_id_0),
    .io_in_id_1(mesh_1_5_io_in_id_1),
    .io_in_last_0(mesh_1_5_io_in_last_0),
    .io_in_last_1(mesh_1_5_io_in_last_1),
    .io_out_a_0(mesh_1_5_io_out_a_0),
    .io_out_a_1(mesh_1_5_io_out_a_1),
    .io_out_c_0(mesh_1_5_io_out_c_0),
    .io_out_c_1(mesh_1_5_io_out_c_1),
    .io_out_b_0(mesh_1_5_io_out_b_0),
    .io_out_b_1(mesh_1_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_5_io_out_control_1_shift),
    .io_out_id_0(mesh_1_5_io_out_id_0),
    .io_out_id_1(mesh_1_5_io_out_id_1),
    .io_out_last_0(mesh_1_5_io_out_last_0),
    .io_out_last_1(mesh_1_5_io_out_last_1),
    .io_in_valid_0(mesh_1_5_io_in_valid_0),
    .io_in_valid_1(mesh_1_5_io_in_valid_1),
    .io_out_valid_0(mesh_1_5_io_out_valid_0),
    .io_out_valid_1(mesh_1_5_io_out_valid_1)
  );
  Tile mesh_1_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_6_clock),
    .io_in_a_0(mesh_1_6_io_in_a_0),
    .io_in_a_1(mesh_1_6_io_in_a_1),
    .io_in_b_0(mesh_1_6_io_in_b_0),
    .io_in_b_1(mesh_1_6_io_in_b_1),
    .io_in_d_0(mesh_1_6_io_in_d_0),
    .io_in_d_1(mesh_1_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_6_io_in_control_1_shift),
    .io_in_id_0(mesh_1_6_io_in_id_0),
    .io_in_id_1(mesh_1_6_io_in_id_1),
    .io_in_last_0(mesh_1_6_io_in_last_0),
    .io_in_last_1(mesh_1_6_io_in_last_1),
    .io_out_a_0(mesh_1_6_io_out_a_0),
    .io_out_a_1(mesh_1_6_io_out_a_1),
    .io_out_c_0(mesh_1_6_io_out_c_0),
    .io_out_c_1(mesh_1_6_io_out_c_1),
    .io_out_b_0(mesh_1_6_io_out_b_0),
    .io_out_b_1(mesh_1_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_6_io_out_control_1_shift),
    .io_out_id_0(mesh_1_6_io_out_id_0),
    .io_out_id_1(mesh_1_6_io_out_id_1),
    .io_out_last_0(mesh_1_6_io_out_last_0),
    .io_out_last_1(mesh_1_6_io_out_last_1),
    .io_in_valid_0(mesh_1_6_io_in_valid_0),
    .io_in_valid_1(mesh_1_6_io_in_valid_1),
    .io_out_valid_0(mesh_1_6_io_out_valid_0),
    .io_out_valid_1(mesh_1_6_io_out_valid_1)
  );
  Tile mesh_1_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_7_clock),
    .io_in_a_0(mesh_1_7_io_in_a_0),
    .io_in_a_1(mesh_1_7_io_in_a_1),
    .io_in_b_0(mesh_1_7_io_in_b_0),
    .io_in_b_1(mesh_1_7_io_in_b_1),
    .io_in_d_0(mesh_1_7_io_in_d_0),
    .io_in_d_1(mesh_1_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_7_io_in_control_1_shift),
    .io_in_id_0(mesh_1_7_io_in_id_0),
    .io_in_id_1(mesh_1_7_io_in_id_1),
    .io_in_last_0(mesh_1_7_io_in_last_0),
    .io_in_last_1(mesh_1_7_io_in_last_1),
    .io_out_a_0(mesh_1_7_io_out_a_0),
    .io_out_a_1(mesh_1_7_io_out_a_1),
    .io_out_c_0(mesh_1_7_io_out_c_0),
    .io_out_c_1(mesh_1_7_io_out_c_1),
    .io_out_b_0(mesh_1_7_io_out_b_0),
    .io_out_b_1(mesh_1_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_7_io_out_control_1_shift),
    .io_out_id_0(mesh_1_7_io_out_id_0),
    .io_out_id_1(mesh_1_7_io_out_id_1),
    .io_out_last_0(mesh_1_7_io_out_last_0),
    .io_out_last_1(mesh_1_7_io_out_last_1),
    .io_in_valid_0(mesh_1_7_io_in_valid_0),
    .io_in_valid_1(mesh_1_7_io_in_valid_1),
    .io_out_valid_0(mesh_1_7_io_out_valid_0),
    .io_out_valid_1(mesh_1_7_io_out_valid_1)
  );
  Tile mesh_1_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_8_clock),
    .io_in_a_0(mesh_1_8_io_in_a_0),
    .io_in_a_1(mesh_1_8_io_in_a_1),
    .io_in_b_0(mesh_1_8_io_in_b_0),
    .io_in_b_1(mesh_1_8_io_in_b_1),
    .io_in_d_0(mesh_1_8_io_in_d_0),
    .io_in_d_1(mesh_1_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_8_io_in_control_1_shift),
    .io_in_id_0(mesh_1_8_io_in_id_0),
    .io_in_id_1(mesh_1_8_io_in_id_1),
    .io_in_last_0(mesh_1_8_io_in_last_0),
    .io_in_last_1(mesh_1_8_io_in_last_1),
    .io_out_a_0(mesh_1_8_io_out_a_0),
    .io_out_a_1(mesh_1_8_io_out_a_1),
    .io_out_c_0(mesh_1_8_io_out_c_0),
    .io_out_c_1(mesh_1_8_io_out_c_1),
    .io_out_b_0(mesh_1_8_io_out_b_0),
    .io_out_b_1(mesh_1_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_8_io_out_control_1_shift),
    .io_out_id_0(mesh_1_8_io_out_id_0),
    .io_out_id_1(mesh_1_8_io_out_id_1),
    .io_out_last_0(mesh_1_8_io_out_last_0),
    .io_out_last_1(mesh_1_8_io_out_last_1),
    .io_in_valid_0(mesh_1_8_io_in_valid_0),
    .io_in_valid_1(mesh_1_8_io_in_valid_1),
    .io_out_valid_0(mesh_1_8_io_out_valid_0),
    .io_out_valid_1(mesh_1_8_io_out_valid_1)
  );
  Tile mesh_1_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_9_clock),
    .io_in_a_0(mesh_1_9_io_in_a_0),
    .io_in_a_1(mesh_1_9_io_in_a_1),
    .io_in_b_0(mesh_1_9_io_in_b_0),
    .io_in_b_1(mesh_1_9_io_in_b_1),
    .io_in_d_0(mesh_1_9_io_in_d_0),
    .io_in_d_1(mesh_1_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_9_io_in_control_1_shift),
    .io_in_id_0(mesh_1_9_io_in_id_0),
    .io_in_id_1(mesh_1_9_io_in_id_1),
    .io_in_last_0(mesh_1_9_io_in_last_0),
    .io_in_last_1(mesh_1_9_io_in_last_1),
    .io_out_a_0(mesh_1_9_io_out_a_0),
    .io_out_a_1(mesh_1_9_io_out_a_1),
    .io_out_c_0(mesh_1_9_io_out_c_0),
    .io_out_c_1(mesh_1_9_io_out_c_1),
    .io_out_b_0(mesh_1_9_io_out_b_0),
    .io_out_b_1(mesh_1_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_9_io_out_control_1_shift),
    .io_out_id_0(mesh_1_9_io_out_id_0),
    .io_out_id_1(mesh_1_9_io_out_id_1),
    .io_out_last_0(mesh_1_9_io_out_last_0),
    .io_out_last_1(mesh_1_9_io_out_last_1),
    .io_in_valid_0(mesh_1_9_io_in_valid_0),
    .io_in_valid_1(mesh_1_9_io_in_valid_1),
    .io_out_valid_0(mesh_1_9_io_out_valid_0),
    .io_out_valid_1(mesh_1_9_io_out_valid_1)
  );
  Tile mesh_1_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_10_clock),
    .io_in_a_0(mesh_1_10_io_in_a_0),
    .io_in_a_1(mesh_1_10_io_in_a_1),
    .io_in_b_0(mesh_1_10_io_in_b_0),
    .io_in_b_1(mesh_1_10_io_in_b_1),
    .io_in_d_0(mesh_1_10_io_in_d_0),
    .io_in_d_1(mesh_1_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_10_io_in_control_1_shift),
    .io_in_id_0(mesh_1_10_io_in_id_0),
    .io_in_id_1(mesh_1_10_io_in_id_1),
    .io_in_last_0(mesh_1_10_io_in_last_0),
    .io_in_last_1(mesh_1_10_io_in_last_1),
    .io_out_a_0(mesh_1_10_io_out_a_0),
    .io_out_a_1(mesh_1_10_io_out_a_1),
    .io_out_c_0(mesh_1_10_io_out_c_0),
    .io_out_c_1(mesh_1_10_io_out_c_1),
    .io_out_b_0(mesh_1_10_io_out_b_0),
    .io_out_b_1(mesh_1_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_10_io_out_control_1_shift),
    .io_out_id_0(mesh_1_10_io_out_id_0),
    .io_out_id_1(mesh_1_10_io_out_id_1),
    .io_out_last_0(mesh_1_10_io_out_last_0),
    .io_out_last_1(mesh_1_10_io_out_last_1),
    .io_in_valid_0(mesh_1_10_io_in_valid_0),
    .io_in_valid_1(mesh_1_10_io_in_valid_1),
    .io_out_valid_0(mesh_1_10_io_out_valid_0),
    .io_out_valid_1(mesh_1_10_io_out_valid_1)
  );
  Tile mesh_1_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_11_clock),
    .io_in_a_0(mesh_1_11_io_in_a_0),
    .io_in_a_1(mesh_1_11_io_in_a_1),
    .io_in_b_0(mesh_1_11_io_in_b_0),
    .io_in_b_1(mesh_1_11_io_in_b_1),
    .io_in_d_0(mesh_1_11_io_in_d_0),
    .io_in_d_1(mesh_1_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_11_io_in_control_1_shift),
    .io_in_id_0(mesh_1_11_io_in_id_0),
    .io_in_id_1(mesh_1_11_io_in_id_1),
    .io_in_last_0(mesh_1_11_io_in_last_0),
    .io_in_last_1(mesh_1_11_io_in_last_1),
    .io_out_a_0(mesh_1_11_io_out_a_0),
    .io_out_a_1(mesh_1_11_io_out_a_1),
    .io_out_c_0(mesh_1_11_io_out_c_0),
    .io_out_c_1(mesh_1_11_io_out_c_1),
    .io_out_b_0(mesh_1_11_io_out_b_0),
    .io_out_b_1(mesh_1_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_11_io_out_control_1_shift),
    .io_out_id_0(mesh_1_11_io_out_id_0),
    .io_out_id_1(mesh_1_11_io_out_id_1),
    .io_out_last_0(mesh_1_11_io_out_last_0),
    .io_out_last_1(mesh_1_11_io_out_last_1),
    .io_in_valid_0(mesh_1_11_io_in_valid_0),
    .io_in_valid_1(mesh_1_11_io_in_valid_1),
    .io_out_valid_0(mesh_1_11_io_out_valid_0),
    .io_out_valid_1(mesh_1_11_io_out_valid_1)
  );
  Tile mesh_1_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_12_clock),
    .io_in_a_0(mesh_1_12_io_in_a_0),
    .io_in_a_1(mesh_1_12_io_in_a_1),
    .io_in_b_0(mesh_1_12_io_in_b_0),
    .io_in_b_1(mesh_1_12_io_in_b_1),
    .io_in_d_0(mesh_1_12_io_in_d_0),
    .io_in_d_1(mesh_1_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_12_io_in_control_1_shift),
    .io_in_id_0(mesh_1_12_io_in_id_0),
    .io_in_id_1(mesh_1_12_io_in_id_1),
    .io_in_last_0(mesh_1_12_io_in_last_0),
    .io_in_last_1(mesh_1_12_io_in_last_1),
    .io_out_a_0(mesh_1_12_io_out_a_0),
    .io_out_a_1(mesh_1_12_io_out_a_1),
    .io_out_c_0(mesh_1_12_io_out_c_0),
    .io_out_c_1(mesh_1_12_io_out_c_1),
    .io_out_b_0(mesh_1_12_io_out_b_0),
    .io_out_b_1(mesh_1_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_12_io_out_control_1_shift),
    .io_out_id_0(mesh_1_12_io_out_id_0),
    .io_out_id_1(mesh_1_12_io_out_id_1),
    .io_out_last_0(mesh_1_12_io_out_last_0),
    .io_out_last_1(mesh_1_12_io_out_last_1),
    .io_in_valid_0(mesh_1_12_io_in_valid_0),
    .io_in_valid_1(mesh_1_12_io_in_valid_1),
    .io_out_valid_0(mesh_1_12_io_out_valid_0),
    .io_out_valid_1(mesh_1_12_io_out_valid_1)
  );
  Tile mesh_1_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_13_clock),
    .io_in_a_0(mesh_1_13_io_in_a_0),
    .io_in_a_1(mesh_1_13_io_in_a_1),
    .io_in_b_0(mesh_1_13_io_in_b_0),
    .io_in_b_1(mesh_1_13_io_in_b_1),
    .io_in_d_0(mesh_1_13_io_in_d_0),
    .io_in_d_1(mesh_1_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_13_io_in_control_1_shift),
    .io_in_id_0(mesh_1_13_io_in_id_0),
    .io_in_id_1(mesh_1_13_io_in_id_1),
    .io_in_last_0(mesh_1_13_io_in_last_0),
    .io_in_last_1(mesh_1_13_io_in_last_1),
    .io_out_a_0(mesh_1_13_io_out_a_0),
    .io_out_a_1(mesh_1_13_io_out_a_1),
    .io_out_c_0(mesh_1_13_io_out_c_0),
    .io_out_c_1(mesh_1_13_io_out_c_1),
    .io_out_b_0(mesh_1_13_io_out_b_0),
    .io_out_b_1(mesh_1_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_13_io_out_control_1_shift),
    .io_out_id_0(mesh_1_13_io_out_id_0),
    .io_out_id_1(mesh_1_13_io_out_id_1),
    .io_out_last_0(mesh_1_13_io_out_last_0),
    .io_out_last_1(mesh_1_13_io_out_last_1),
    .io_in_valid_0(mesh_1_13_io_in_valid_0),
    .io_in_valid_1(mesh_1_13_io_in_valid_1),
    .io_out_valid_0(mesh_1_13_io_out_valid_0),
    .io_out_valid_1(mesh_1_13_io_out_valid_1)
  );
  Tile mesh_1_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_14_clock),
    .io_in_a_0(mesh_1_14_io_in_a_0),
    .io_in_a_1(mesh_1_14_io_in_a_1),
    .io_in_b_0(mesh_1_14_io_in_b_0),
    .io_in_b_1(mesh_1_14_io_in_b_1),
    .io_in_d_0(mesh_1_14_io_in_d_0),
    .io_in_d_1(mesh_1_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_14_io_in_control_1_shift),
    .io_in_id_0(mesh_1_14_io_in_id_0),
    .io_in_id_1(mesh_1_14_io_in_id_1),
    .io_in_last_0(mesh_1_14_io_in_last_0),
    .io_in_last_1(mesh_1_14_io_in_last_1),
    .io_out_a_0(mesh_1_14_io_out_a_0),
    .io_out_a_1(mesh_1_14_io_out_a_1),
    .io_out_c_0(mesh_1_14_io_out_c_0),
    .io_out_c_1(mesh_1_14_io_out_c_1),
    .io_out_b_0(mesh_1_14_io_out_b_0),
    .io_out_b_1(mesh_1_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_14_io_out_control_1_shift),
    .io_out_id_0(mesh_1_14_io_out_id_0),
    .io_out_id_1(mesh_1_14_io_out_id_1),
    .io_out_last_0(mesh_1_14_io_out_last_0),
    .io_out_last_1(mesh_1_14_io_out_last_1),
    .io_in_valid_0(mesh_1_14_io_in_valid_0),
    .io_in_valid_1(mesh_1_14_io_in_valid_1),
    .io_out_valid_0(mesh_1_14_io_out_valid_0),
    .io_out_valid_1(mesh_1_14_io_out_valid_1)
  );
  Tile mesh_1_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_1_15_clock),
    .io_in_a_0(mesh_1_15_io_in_a_0),
    .io_in_a_1(mesh_1_15_io_in_a_1),
    .io_in_b_0(mesh_1_15_io_in_b_0),
    .io_in_b_1(mesh_1_15_io_in_b_1),
    .io_in_d_0(mesh_1_15_io_in_d_0),
    .io_in_d_1(mesh_1_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_15_io_in_control_1_shift),
    .io_in_id_0(mesh_1_15_io_in_id_0),
    .io_in_id_1(mesh_1_15_io_in_id_1),
    .io_in_last_0(mesh_1_15_io_in_last_0),
    .io_in_last_1(mesh_1_15_io_in_last_1),
    .io_out_a_0(mesh_1_15_io_out_a_0),
    .io_out_a_1(mesh_1_15_io_out_a_1),
    .io_out_c_0(mesh_1_15_io_out_c_0),
    .io_out_c_1(mesh_1_15_io_out_c_1),
    .io_out_b_0(mesh_1_15_io_out_b_0),
    .io_out_b_1(mesh_1_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_15_io_out_control_1_shift),
    .io_out_id_0(mesh_1_15_io_out_id_0),
    .io_out_id_1(mesh_1_15_io_out_id_1),
    .io_out_last_0(mesh_1_15_io_out_last_0),
    .io_out_last_1(mesh_1_15_io_out_last_1),
    .io_in_valid_0(mesh_1_15_io_in_valid_0),
    .io_in_valid_1(mesh_1_15_io_in_valid_1),
    .io_out_valid_0(mesh_1_15_io_out_valid_0),
    .io_out_valid_1(mesh_1_15_io_out_valid_1)
  );
  Tile mesh_2_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_0_clock),
    .io_in_a_0(mesh_2_0_io_in_a_0),
    .io_in_a_1(mesh_2_0_io_in_a_1),
    .io_in_b_0(mesh_2_0_io_in_b_0),
    .io_in_b_1(mesh_2_0_io_in_b_1),
    .io_in_d_0(mesh_2_0_io_in_d_0),
    .io_in_d_1(mesh_2_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_0_io_in_control_1_shift),
    .io_in_id_0(mesh_2_0_io_in_id_0),
    .io_in_id_1(mesh_2_0_io_in_id_1),
    .io_in_last_0(mesh_2_0_io_in_last_0),
    .io_in_last_1(mesh_2_0_io_in_last_1),
    .io_out_a_0(mesh_2_0_io_out_a_0),
    .io_out_a_1(mesh_2_0_io_out_a_1),
    .io_out_c_0(mesh_2_0_io_out_c_0),
    .io_out_c_1(mesh_2_0_io_out_c_1),
    .io_out_b_0(mesh_2_0_io_out_b_0),
    .io_out_b_1(mesh_2_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_0_io_out_control_1_shift),
    .io_out_id_0(mesh_2_0_io_out_id_0),
    .io_out_id_1(mesh_2_0_io_out_id_1),
    .io_out_last_0(mesh_2_0_io_out_last_0),
    .io_out_last_1(mesh_2_0_io_out_last_1),
    .io_in_valid_0(mesh_2_0_io_in_valid_0),
    .io_in_valid_1(mesh_2_0_io_in_valid_1),
    .io_out_valid_0(mesh_2_0_io_out_valid_0),
    .io_out_valid_1(mesh_2_0_io_out_valid_1)
  );
  Tile mesh_2_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_1_clock),
    .io_in_a_0(mesh_2_1_io_in_a_0),
    .io_in_a_1(mesh_2_1_io_in_a_1),
    .io_in_b_0(mesh_2_1_io_in_b_0),
    .io_in_b_1(mesh_2_1_io_in_b_1),
    .io_in_d_0(mesh_2_1_io_in_d_0),
    .io_in_d_1(mesh_2_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_1_io_in_control_1_shift),
    .io_in_id_0(mesh_2_1_io_in_id_0),
    .io_in_id_1(mesh_2_1_io_in_id_1),
    .io_in_last_0(mesh_2_1_io_in_last_0),
    .io_in_last_1(mesh_2_1_io_in_last_1),
    .io_out_a_0(mesh_2_1_io_out_a_0),
    .io_out_a_1(mesh_2_1_io_out_a_1),
    .io_out_c_0(mesh_2_1_io_out_c_0),
    .io_out_c_1(mesh_2_1_io_out_c_1),
    .io_out_b_0(mesh_2_1_io_out_b_0),
    .io_out_b_1(mesh_2_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_1_io_out_control_1_shift),
    .io_out_id_0(mesh_2_1_io_out_id_0),
    .io_out_id_1(mesh_2_1_io_out_id_1),
    .io_out_last_0(mesh_2_1_io_out_last_0),
    .io_out_last_1(mesh_2_1_io_out_last_1),
    .io_in_valid_0(mesh_2_1_io_in_valid_0),
    .io_in_valid_1(mesh_2_1_io_in_valid_1),
    .io_out_valid_0(mesh_2_1_io_out_valid_0),
    .io_out_valid_1(mesh_2_1_io_out_valid_1)
  );
  Tile mesh_2_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_2_clock),
    .io_in_a_0(mesh_2_2_io_in_a_0),
    .io_in_a_1(mesh_2_2_io_in_a_1),
    .io_in_b_0(mesh_2_2_io_in_b_0),
    .io_in_b_1(mesh_2_2_io_in_b_1),
    .io_in_d_0(mesh_2_2_io_in_d_0),
    .io_in_d_1(mesh_2_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_2_io_in_control_1_shift),
    .io_in_id_0(mesh_2_2_io_in_id_0),
    .io_in_id_1(mesh_2_2_io_in_id_1),
    .io_in_last_0(mesh_2_2_io_in_last_0),
    .io_in_last_1(mesh_2_2_io_in_last_1),
    .io_out_a_0(mesh_2_2_io_out_a_0),
    .io_out_a_1(mesh_2_2_io_out_a_1),
    .io_out_c_0(mesh_2_2_io_out_c_0),
    .io_out_c_1(mesh_2_2_io_out_c_1),
    .io_out_b_0(mesh_2_2_io_out_b_0),
    .io_out_b_1(mesh_2_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_2_io_out_control_1_shift),
    .io_out_id_0(mesh_2_2_io_out_id_0),
    .io_out_id_1(mesh_2_2_io_out_id_1),
    .io_out_last_0(mesh_2_2_io_out_last_0),
    .io_out_last_1(mesh_2_2_io_out_last_1),
    .io_in_valid_0(mesh_2_2_io_in_valid_0),
    .io_in_valid_1(mesh_2_2_io_in_valid_1),
    .io_out_valid_0(mesh_2_2_io_out_valid_0),
    .io_out_valid_1(mesh_2_2_io_out_valid_1)
  );
  Tile mesh_2_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_3_clock),
    .io_in_a_0(mesh_2_3_io_in_a_0),
    .io_in_a_1(mesh_2_3_io_in_a_1),
    .io_in_b_0(mesh_2_3_io_in_b_0),
    .io_in_b_1(mesh_2_3_io_in_b_1),
    .io_in_d_0(mesh_2_3_io_in_d_0),
    .io_in_d_1(mesh_2_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_3_io_in_control_1_shift),
    .io_in_id_0(mesh_2_3_io_in_id_0),
    .io_in_id_1(mesh_2_3_io_in_id_1),
    .io_in_last_0(mesh_2_3_io_in_last_0),
    .io_in_last_1(mesh_2_3_io_in_last_1),
    .io_out_a_0(mesh_2_3_io_out_a_0),
    .io_out_a_1(mesh_2_3_io_out_a_1),
    .io_out_c_0(mesh_2_3_io_out_c_0),
    .io_out_c_1(mesh_2_3_io_out_c_1),
    .io_out_b_0(mesh_2_3_io_out_b_0),
    .io_out_b_1(mesh_2_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_3_io_out_control_1_shift),
    .io_out_id_0(mesh_2_3_io_out_id_0),
    .io_out_id_1(mesh_2_3_io_out_id_1),
    .io_out_last_0(mesh_2_3_io_out_last_0),
    .io_out_last_1(mesh_2_3_io_out_last_1),
    .io_in_valid_0(mesh_2_3_io_in_valid_0),
    .io_in_valid_1(mesh_2_3_io_in_valid_1),
    .io_out_valid_0(mesh_2_3_io_out_valid_0),
    .io_out_valid_1(mesh_2_3_io_out_valid_1)
  );
  Tile mesh_2_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_4_clock),
    .io_in_a_0(mesh_2_4_io_in_a_0),
    .io_in_a_1(mesh_2_4_io_in_a_1),
    .io_in_b_0(mesh_2_4_io_in_b_0),
    .io_in_b_1(mesh_2_4_io_in_b_1),
    .io_in_d_0(mesh_2_4_io_in_d_0),
    .io_in_d_1(mesh_2_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_4_io_in_control_1_shift),
    .io_in_id_0(mesh_2_4_io_in_id_0),
    .io_in_id_1(mesh_2_4_io_in_id_1),
    .io_in_last_0(mesh_2_4_io_in_last_0),
    .io_in_last_1(mesh_2_4_io_in_last_1),
    .io_out_a_0(mesh_2_4_io_out_a_0),
    .io_out_a_1(mesh_2_4_io_out_a_1),
    .io_out_c_0(mesh_2_4_io_out_c_0),
    .io_out_c_1(mesh_2_4_io_out_c_1),
    .io_out_b_0(mesh_2_4_io_out_b_0),
    .io_out_b_1(mesh_2_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_4_io_out_control_1_shift),
    .io_out_id_0(mesh_2_4_io_out_id_0),
    .io_out_id_1(mesh_2_4_io_out_id_1),
    .io_out_last_0(mesh_2_4_io_out_last_0),
    .io_out_last_1(mesh_2_4_io_out_last_1),
    .io_in_valid_0(mesh_2_4_io_in_valid_0),
    .io_in_valid_1(mesh_2_4_io_in_valid_1),
    .io_out_valid_0(mesh_2_4_io_out_valid_0),
    .io_out_valid_1(mesh_2_4_io_out_valid_1)
  );
  Tile mesh_2_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_5_clock),
    .io_in_a_0(mesh_2_5_io_in_a_0),
    .io_in_a_1(mesh_2_5_io_in_a_1),
    .io_in_b_0(mesh_2_5_io_in_b_0),
    .io_in_b_1(mesh_2_5_io_in_b_1),
    .io_in_d_0(mesh_2_5_io_in_d_0),
    .io_in_d_1(mesh_2_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_5_io_in_control_1_shift),
    .io_in_id_0(mesh_2_5_io_in_id_0),
    .io_in_id_1(mesh_2_5_io_in_id_1),
    .io_in_last_0(mesh_2_5_io_in_last_0),
    .io_in_last_1(mesh_2_5_io_in_last_1),
    .io_out_a_0(mesh_2_5_io_out_a_0),
    .io_out_a_1(mesh_2_5_io_out_a_1),
    .io_out_c_0(mesh_2_5_io_out_c_0),
    .io_out_c_1(mesh_2_5_io_out_c_1),
    .io_out_b_0(mesh_2_5_io_out_b_0),
    .io_out_b_1(mesh_2_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_5_io_out_control_1_shift),
    .io_out_id_0(mesh_2_5_io_out_id_0),
    .io_out_id_1(mesh_2_5_io_out_id_1),
    .io_out_last_0(mesh_2_5_io_out_last_0),
    .io_out_last_1(mesh_2_5_io_out_last_1),
    .io_in_valid_0(mesh_2_5_io_in_valid_0),
    .io_in_valid_1(mesh_2_5_io_in_valid_1),
    .io_out_valid_0(mesh_2_5_io_out_valid_0),
    .io_out_valid_1(mesh_2_5_io_out_valid_1)
  );
  Tile mesh_2_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_6_clock),
    .io_in_a_0(mesh_2_6_io_in_a_0),
    .io_in_a_1(mesh_2_6_io_in_a_1),
    .io_in_b_0(mesh_2_6_io_in_b_0),
    .io_in_b_1(mesh_2_6_io_in_b_1),
    .io_in_d_0(mesh_2_6_io_in_d_0),
    .io_in_d_1(mesh_2_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_6_io_in_control_1_shift),
    .io_in_id_0(mesh_2_6_io_in_id_0),
    .io_in_id_1(mesh_2_6_io_in_id_1),
    .io_in_last_0(mesh_2_6_io_in_last_0),
    .io_in_last_1(mesh_2_6_io_in_last_1),
    .io_out_a_0(mesh_2_6_io_out_a_0),
    .io_out_a_1(mesh_2_6_io_out_a_1),
    .io_out_c_0(mesh_2_6_io_out_c_0),
    .io_out_c_1(mesh_2_6_io_out_c_1),
    .io_out_b_0(mesh_2_6_io_out_b_0),
    .io_out_b_1(mesh_2_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_6_io_out_control_1_shift),
    .io_out_id_0(mesh_2_6_io_out_id_0),
    .io_out_id_1(mesh_2_6_io_out_id_1),
    .io_out_last_0(mesh_2_6_io_out_last_0),
    .io_out_last_1(mesh_2_6_io_out_last_1),
    .io_in_valid_0(mesh_2_6_io_in_valid_0),
    .io_in_valid_1(mesh_2_6_io_in_valid_1),
    .io_out_valid_0(mesh_2_6_io_out_valid_0),
    .io_out_valid_1(mesh_2_6_io_out_valid_1)
  );
  Tile mesh_2_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_7_clock),
    .io_in_a_0(mesh_2_7_io_in_a_0),
    .io_in_a_1(mesh_2_7_io_in_a_1),
    .io_in_b_0(mesh_2_7_io_in_b_0),
    .io_in_b_1(mesh_2_7_io_in_b_1),
    .io_in_d_0(mesh_2_7_io_in_d_0),
    .io_in_d_1(mesh_2_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_7_io_in_control_1_shift),
    .io_in_id_0(mesh_2_7_io_in_id_0),
    .io_in_id_1(mesh_2_7_io_in_id_1),
    .io_in_last_0(mesh_2_7_io_in_last_0),
    .io_in_last_1(mesh_2_7_io_in_last_1),
    .io_out_a_0(mesh_2_7_io_out_a_0),
    .io_out_a_1(mesh_2_7_io_out_a_1),
    .io_out_c_0(mesh_2_7_io_out_c_0),
    .io_out_c_1(mesh_2_7_io_out_c_1),
    .io_out_b_0(mesh_2_7_io_out_b_0),
    .io_out_b_1(mesh_2_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_7_io_out_control_1_shift),
    .io_out_id_0(mesh_2_7_io_out_id_0),
    .io_out_id_1(mesh_2_7_io_out_id_1),
    .io_out_last_0(mesh_2_7_io_out_last_0),
    .io_out_last_1(mesh_2_7_io_out_last_1),
    .io_in_valid_0(mesh_2_7_io_in_valid_0),
    .io_in_valid_1(mesh_2_7_io_in_valid_1),
    .io_out_valid_0(mesh_2_7_io_out_valid_0),
    .io_out_valid_1(mesh_2_7_io_out_valid_1)
  );
  Tile mesh_2_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_8_clock),
    .io_in_a_0(mesh_2_8_io_in_a_0),
    .io_in_a_1(mesh_2_8_io_in_a_1),
    .io_in_b_0(mesh_2_8_io_in_b_0),
    .io_in_b_1(mesh_2_8_io_in_b_1),
    .io_in_d_0(mesh_2_8_io_in_d_0),
    .io_in_d_1(mesh_2_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_8_io_in_control_1_shift),
    .io_in_id_0(mesh_2_8_io_in_id_0),
    .io_in_id_1(mesh_2_8_io_in_id_1),
    .io_in_last_0(mesh_2_8_io_in_last_0),
    .io_in_last_1(mesh_2_8_io_in_last_1),
    .io_out_a_0(mesh_2_8_io_out_a_0),
    .io_out_a_1(mesh_2_8_io_out_a_1),
    .io_out_c_0(mesh_2_8_io_out_c_0),
    .io_out_c_1(mesh_2_8_io_out_c_1),
    .io_out_b_0(mesh_2_8_io_out_b_0),
    .io_out_b_1(mesh_2_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_8_io_out_control_1_shift),
    .io_out_id_0(mesh_2_8_io_out_id_0),
    .io_out_id_1(mesh_2_8_io_out_id_1),
    .io_out_last_0(mesh_2_8_io_out_last_0),
    .io_out_last_1(mesh_2_8_io_out_last_1),
    .io_in_valid_0(mesh_2_8_io_in_valid_0),
    .io_in_valid_1(mesh_2_8_io_in_valid_1),
    .io_out_valid_0(mesh_2_8_io_out_valid_0),
    .io_out_valid_1(mesh_2_8_io_out_valid_1)
  );
  Tile mesh_2_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_9_clock),
    .io_in_a_0(mesh_2_9_io_in_a_0),
    .io_in_a_1(mesh_2_9_io_in_a_1),
    .io_in_b_0(mesh_2_9_io_in_b_0),
    .io_in_b_1(mesh_2_9_io_in_b_1),
    .io_in_d_0(mesh_2_9_io_in_d_0),
    .io_in_d_1(mesh_2_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_9_io_in_control_1_shift),
    .io_in_id_0(mesh_2_9_io_in_id_0),
    .io_in_id_1(mesh_2_9_io_in_id_1),
    .io_in_last_0(mesh_2_9_io_in_last_0),
    .io_in_last_1(mesh_2_9_io_in_last_1),
    .io_out_a_0(mesh_2_9_io_out_a_0),
    .io_out_a_1(mesh_2_9_io_out_a_1),
    .io_out_c_0(mesh_2_9_io_out_c_0),
    .io_out_c_1(mesh_2_9_io_out_c_1),
    .io_out_b_0(mesh_2_9_io_out_b_0),
    .io_out_b_1(mesh_2_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_9_io_out_control_1_shift),
    .io_out_id_0(mesh_2_9_io_out_id_0),
    .io_out_id_1(mesh_2_9_io_out_id_1),
    .io_out_last_0(mesh_2_9_io_out_last_0),
    .io_out_last_1(mesh_2_9_io_out_last_1),
    .io_in_valid_0(mesh_2_9_io_in_valid_0),
    .io_in_valid_1(mesh_2_9_io_in_valid_1),
    .io_out_valid_0(mesh_2_9_io_out_valid_0),
    .io_out_valid_1(mesh_2_9_io_out_valid_1)
  );
  Tile mesh_2_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_10_clock),
    .io_in_a_0(mesh_2_10_io_in_a_0),
    .io_in_a_1(mesh_2_10_io_in_a_1),
    .io_in_b_0(mesh_2_10_io_in_b_0),
    .io_in_b_1(mesh_2_10_io_in_b_1),
    .io_in_d_0(mesh_2_10_io_in_d_0),
    .io_in_d_1(mesh_2_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_10_io_in_control_1_shift),
    .io_in_id_0(mesh_2_10_io_in_id_0),
    .io_in_id_1(mesh_2_10_io_in_id_1),
    .io_in_last_0(mesh_2_10_io_in_last_0),
    .io_in_last_1(mesh_2_10_io_in_last_1),
    .io_out_a_0(mesh_2_10_io_out_a_0),
    .io_out_a_1(mesh_2_10_io_out_a_1),
    .io_out_c_0(mesh_2_10_io_out_c_0),
    .io_out_c_1(mesh_2_10_io_out_c_1),
    .io_out_b_0(mesh_2_10_io_out_b_0),
    .io_out_b_1(mesh_2_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_10_io_out_control_1_shift),
    .io_out_id_0(mesh_2_10_io_out_id_0),
    .io_out_id_1(mesh_2_10_io_out_id_1),
    .io_out_last_0(mesh_2_10_io_out_last_0),
    .io_out_last_1(mesh_2_10_io_out_last_1),
    .io_in_valid_0(mesh_2_10_io_in_valid_0),
    .io_in_valid_1(mesh_2_10_io_in_valid_1),
    .io_out_valid_0(mesh_2_10_io_out_valid_0),
    .io_out_valid_1(mesh_2_10_io_out_valid_1)
  );
  Tile mesh_2_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_11_clock),
    .io_in_a_0(mesh_2_11_io_in_a_0),
    .io_in_a_1(mesh_2_11_io_in_a_1),
    .io_in_b_0(mesh_2_11_io_in_b_0),
    .io_in_b_1(mesh_2_11_io_in_b_1),
    .io_in_d_0(mesh_2_11_io_in_d_0),
    .io_in_d_1(mesh_2_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_11_io_in_control_1_shift),
    .io_in_id_0(mesh_2_11_io_in_id_0),
    .io_in_id_1(mesh_2_11_io_in_id_1),
    .io_in_last_0(mesh_2_11_io_in_last_0),
    .io_in_last_1(mesh_2_11_io_in_last_1),
    .io_out_a_0(mesh_2_11_io_out_a_0),
    .io_out_a_1(mesh_2_11_io_out_a_1),
    .io_out_c_0(mesh_2_11_io_out_c_0),
    .io_out_c_1(mesh_2_11_io_out_c_1),
    .io_out_b_0(mesh_2_11_io_out_b_0),
    .io_out_b_1(mesh_2_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_11_io_out_control_1_shift),
    .io_out_id_0(mesh_2_11_io_out_id_0),
    .io_out_id_1(mesh_2_11_io_out_id_1),
    .io_out_last_0(mesh_2_11_io_out_last_0),
    .io_out_last_1(mesh_2_11_io_out_last_1),
    .io_in_valid_0(mesh_2_11_io_in_valid_0),
    .io_in_valid_1(mesh_2_11_io_in_valid_1),
    .io_out_valid_0(mesh_2_11_io_out_valid_0),
    .io_out_valid_1(mesh_2_11_io_out_valid_1)
  );
  Tile mesh_2_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_12_clock),
    .io_in_a_0(mesh_2_12_io_in_a_0),
    .io_in_a_1(mesh_2_12_io_in_a_1),
    .io_in_b_0(mesh_2_12_io_in_b_0),
    .io_in_b_1(mesh_2_12_io_in_b_1),
    .io_in_d_0(mesh_2_12_io_in_d_0),
    .io_in_d_1(mesh_2_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_12_io_in_control_1_shift),
    .io_in_id_0(mesh_2_12_io_in_id_0),
    .io_in_id_1(mesh_2_12_io_in_id_1),
    .io_in_last_0(mesh_2_12_io_in_last_0),
    .io_in_last_1(mesh_2_12_io_in_last_1),
    .io_out_a_0(mesh_2_12_io_out_a_0),
    .io_out_a_1(mesh_2_12_io_out_a_1),
    .io_out_c_0(mesh_2_12_io_out_c_0),
    .io_out_c_1(mesh_2_12_io_out_c_1),
    .io_out_b_0(mesh_2_12_io_out_b_0),
    .io_out_b_1(mesh_2_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_12_io_out_control_1_shift),
    .io_out_id_0(mesh_2_12_io_out_id_0),
    .io_out_id_1(mesh_2_12_io_out_id_1),
    .io_out_last_0(mesh_2_12_io_out_last_0),
    .io_out_last_1(mesh_2_12_io_out_last_1),
    .io_in_valid_0(mesh_2_12_io_in_valid_0),
    .io_in_valid_1(mesh_2_12_io_in_valid_1),
    .io_out_valid_0(mesh_2_12_io_out_valid_0),
    .io_out_valid_1(mesh_2_12_io_out_valid_1)
  );
  Tile mesh_2_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_13_clock),
    .io_in_a_0(mesh_2_13_io_in_a_0),
    .io_in_a_1(mesh_2_13_io_in_a_1),
    .io_in_b_0(mesh_2_13_io_in_b_0),
    .io_in_b_1(mesh_2_13_io_in_b_1),
    .io_in_d_0(mesh_2_13_io_in_d_0),
    .io_in_d_1(mesh_2_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_13_io_in_control_1_shift),
    .io_in_id_0(mesh_2_13_io_in_id_0),
    .io_in_id_1(mesh_2_13_io_in_id_1),
    .io_in_last_0(mesh_2_13_io_in_last_0),
    .io_in_last_1(mesh_2_13_io_in_last_1),
    .io_out_a_0(mesh_2_13_io_out_a_0),
    .io_out_a_1(mesh_2_13_io_out_a_1),
    .io_out_c_0(mesh_2_13_io_out_c_0),
    .io_out_c_1(mesh_2_13_io_out_c_1),
    .io_out_b_0(mesh_2_13_io_out_b_0),
    .io_out_b_1(mesh_2_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_13_io_out_control_1_shift),
    .io_out_id_0(mesh_2_13_io_out_id_0),
    .io_out_id_1(mesh_2_13_io_out_id_1),
    .io_out_last_0(mesh_2_13_io_out_last_0),
    .io_out_last_1(mesh_2_13_io_out_last_1),
    .io_in_valid_0(mesh_2_13_io_in_valid_0),
    .io_in_valid_1(mesh_2_13_io_in_valid_1),
    .io_out_valid_0(mesh_2_13_io_out_valid_0),
    .io_out_valid_1(mesh_2_13_io_out_valid_1)
  );
  Tile mesh_2_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_14_clock),
    .io_in_a_0(mesh_2_14_io_in_a_0),
    .io_in_a_1(mesh_2_14_io_in_a_1),
    .io_in_b_0(mesh_2_14_io_in_b_0),
    .io_in_b_1(mesh_2_14_io_in_b_1),
    .io_in_d_0(mesh_2_14_io_in_d_0),
    .io_in_d_1(mesh_2_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_14_io_in_control_1_shift),
    .io_in_id_0(mesh_2_14_io_in_id_0),
    .io_in_id_1(mesh_2_14_io_in_id_1),
    .io_in_last_0(mesh_2_14_io_in_last_0),
    .io_in_last_1(mesh_2_14_io_in_last_1),
    .io_out_a_0(mesh_2_14_io_out_a_0),
    .io_out_a_1(mesh_2_14_io_out_a_1),
    .io_out_c_0(mesh_2_14_io_out_c_0),
    .io_out_c_1(mesh_2_14_io_out_c_1),
    .io_out_b_0(mesh_2_14_io_out_b_0),
    .io_out_b_1(mesh_2_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_14_io_out_control_1_shift),
    .io_out_id_0(mesh_2_14_io_out_id_0),
    .io_out_id_1(mesh_2_14_io_out_id_1),
    .io_out_last_0(mesh_2_14_io_out_last_0),
    .io_out_last_1(mesh_2_14_io_out_last_1),
    .io_in_valid_0(mesh_2_14_io_in_valid_0),
    .io_in_valid_1(mesh_2_14_io_in_valid_1),
    .io_out_valid_0(mesh_2_14_io_out_valid_0),
    .io_out_valid_1(mesh_2_14_io_out_valid_1)
  );
  Tile mesh_2_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_2_15_clock),
    .io_in_a_0(mesh_2_15_io_in_a_0),
    .io_in_a_1(mesh_2_15_io_in_a_1),
    .io_in_b_0(mesh_2_15_io_in_b_0),
    .io_in_b_1(mesh_2_15_io_in_b_1),
    .io_in_d_0(mesh_2_15_io_in_d_0),
    .io_in_d_1(mesh_2_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_2_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_2_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_2_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_2_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_2_15_io_in_control_1_shift),
    .io_in_id_0(mesh_2_15_io_in_id_0),
    .io_in_id_1(mesh_2_15_io_in_id_1),
    .io_in_last_0(mesh_2_15_io_in_last_0),
    .io_in_last_1(mesh_2_15_io_in_last_1),
    .io_out_a_0(mesh_2_15_io_out_a_0),
    .io_out_a_1(mesh_2_15_io_out_a_1),
    .io_out_c_0(mesh_2_15_io_out_c_0),
    .io_out_c_1(mesh_2_15_io_out_c_1),
    .io_out_b_0(mesh_2_15_io_out_b_0),
    .io_out_b_1(mesh_2_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_2_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_2_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_2_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_2_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_2_15_io_out_control_1_shift),
    .io_out_id_0(mesh_2_15_io_out_id_0),
    .io_out_id_1(mesh_2_15_io_out_id_1),
    .io_out_last_0(mesh_2_15_io_out_last_0),
    .io_out_last_1(mesh_2_15_io_out_last_1),
    .io_in_valid_0(mesh_2_15_io_in_valid_0),
    .io_in_valid_1(mesh_2_15_io_in_valid_1),
    .io_out_valid_0(mesh_2_15_io_out_valid_0),
    .io_out_valid_1(mesh_2_15_io_out_valid_1)
  );
  Tile mesh_3_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_0_clock),
    .io_in_a_0(mesh_3_0_io_in_a_0),
    .io_in_a_1(mesh_3_0_io_in_a_1),
    .io_in_b_0(mesh_3_0_io_in_b_0),
    .io_in_b_1(mesh_3_0_io_in_b_1),
    .io_in_d_0(mesh_3_0_io_in_d_0),
    .io_in_d_1(mesh_3_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_0_io_in_control_1_shift),
    .io_in_id_0(mesh_3_0_io_in_id_0),
    .io_in_id_1(mesh_3_0_io_in_id_1),
    .io_in_last_0(mesh_3_0_io_in_last_0),
    .io_in_last_1(mesh_3_0_io_in_last_1),
    .io_out_a_0(mesh_3_0_io_out_a_0),
    .io_out_a_1(mesh_3_0_io_out_a_1),
    .io_out_c_0(mesh_3_0_io_out_c_0),
    .io_out_c_1(mesh_3_0_io_out_c_1),
    .io_out_b_0(mesh_3_0_io_out_b_0),
    .io_out_b_1(mesh_3_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_0_io_out_control_1_shift),
    .io_out_id_0(mesh_3_0_io_out_id_0),
    .io_out_id_1(mesh_3_0_io_out_id_1),
    .io_out_last_0(mesh_3_0_io_out_last_0),
    .io_out_last_1(mesh_3_0_io_out_last_1),
    .io_in_valid_0(mesh_3_0_io_in_valid_0),
    .io_in_valid_1(mesh_3_0_io_in_valid_1),
    .io_out_valid_0(mesh_3_0_io_out_valid_0),
    .io_out_valid_1(mesh_3_0_io_out_valid_1)
  );
  Tile mesh_3_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_1_clock),
    .io_in_a_0(mesh_3_1_io_in_a_0),
    .io_in_a_1(mesh_3_1_io_in_a_1),
    .io_in_b_0(mesh_3_1_io_in_b_0),
    .io_in_b_1(mesh_3_1_io_in_b_1),
    .io_in_d_0(mesh_3_1_io_in_d_0),
    .io_in_d_1(mesh_3_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_1_io_in_control_1_shift),
    .io_in_id_0(mesh_3_1_io_in_id_0),
    .io_in_id_1(mesh_3_1_io_in_id_1),
    .io_in_last_0(mesh_3_1_io_in_last_0),
    .io_in_last_1(mesh_3_1_io_in_last_1),
    .io_out_a_0(mesh_3_1_io_out_a_0),
    .io_out_a_1(mesh_3_1_io_out_a_1),
    .io_out_c_0(mesh_3_1_io_out_c_0),
    .io_out_c_1(mesh_3_1_io_out_c_1),
    .io_out_b_0(mesh_3_1_io_out_b_0),
    .io_out_b_1(mesh_3_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_1_io_out_control_1_shift),
    .io_out_id_0(mesh_3_1_io_out_id_0),
    .io_out_id_1(mesh_3_1_io_out_id_1),
    .io_out_last_0(mesh_3_1_io_out_last_0),
    .io_out_last_1(mesh_3_1_io_out_last_1),
    .io_in_valid_0(mesh_3_1_io_in_valid_0),
    .io_in_valid_1(mesh_3_1_io_in_valid_1),
    .io_out_valid_0(mesh_3_1_io_out_valid_0),
    .io_out_valid_1(mesh_3_1_io_out_valid_1)
  );
  Tile mesh_3_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_2_clock),
    .io_in_a_0(mesh_3_2_io_in_a_0),
    .io_in_a_1(mesh_3_2_io_in_a_1),
    .io_in_b_0(mesh_3_2_io_in_b_0),
    .io_in_b_1(mesh_3_2_io_in_b_1),
    .io_in_d_0(mesh_3_2_io_in_d_0),
    .io_in_d_1(mesh_3_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_2_io_in_control_1_shift),
    .io_in_id_0(mesh_3_2_io_in_id_0),
    .io_in_id_1(mesh_3_2_io_in_id_1),
    .io_in_last_0(mesh_3_2_io_in_last_0),
    .io_in_last_1(mesh_3_2_io_in_last_1),
    .io_out_a_0(mesh_3_2_io_out_a_0),
    .io_out_a_1(mesh_3_2_io_out_a_1),
    .io_out_c_0(mesh_3_2_io_out_c_0),
    .io_out_c_1(mesh_3_2_io_out_c_1),
    .io_out_b_0(mesh_3_2_io_out_b_0),
    .io_out_b_1(mesh_3_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_2_io_out_control_1_shift),
    .io_out_id_0(mesh_3_2_io_out_id_0),
    .io_out_id_1(mesh_3_2_io_out_id_1),
    .io_out_last_0(mesh_3_2_io_out_last_0),
    .io_out_last_1(mesh_3_2_io_out_last_1),
    .io_in_valid_0(mesh_3_2_io_in_valid_0),
    .io_in_valid_1(mesh_3_2_io_in_valid_1),
    .io_out_valid_0(mesh_3_2_io_out_valid_0),
    .io_out_valid_1(mesh_3_2_io_out_valid_1)
  );
  Tile mesh_3_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_3_clock),
    .io_in_a_0(mesh_3_3_io_in_a_0),
    .io_in_a_1(mesh_3_3_io_in_a_1),
    .io_in_b_0(mesh_3_3_io_in_b_0),
    .io_in_b_1(mesh_3_3_io_in_b_1),
    .io_in_d_0(mesh_3_3_io_in_d_0),
    .io_in_d_1(mesh_3_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_3_io_in_control_1_shift),
    .io_in_id_0(mesh_3_3_io_in_id_0),
    .io_in_id_1(mesh_3_3_io_in_id_1),
    .io_in_last_0(mesh_3_3_io_in_last_0),
    .io_in_last_1(mesh_3_3_io_in_last_1),
    .io_out_a_0(mesh_3_3_io_out_a_0),
    .io_out_a_1(mesh_3_3_io_out_a_1),
    .io_out_c_0(mesh_3_3_io_out_c_0),
    .io_out_c_1(mesh_3_3_io_out_c_1),
    .io_out_b_0(mesh_3_3_io_out_b_0),
    .io_out_b_1(mesh_3_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_3_io_out_control_1_shift),
    .io_out_id_0(mesh_3_3_io_out_id_0),
    .io_out_id_1(mesh_3_3_io_out_id_1),
    .io_out_last_0(mesh_3_3_io_out_last_0),
    .io_out_last_1(mesh_3_3_io_out_last_1),
    .io_in_valid_0(mesh_3_3_io_in_valid_0),
    .io_in_valid_1(mesh_3_3_io_in_valid_1),
    .io_out_valid_0(mesh_3_3_io_out_valid_0),
    .io_out_valid_1(mesh_3_3_io_out_valid_1)
  );
  Tile mesh_3_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_4_clock),
    .io_in_a_0(mesh_3_4_io_in_a_0),
    .io_in_a_1(mesh_3_4_io_in_a_1),
    .io_in_b_0(mesh_3_4_io_in_b_0),
    .io_in_b_1(mesh_3_4_io_in_b_1),
    .io_in_d_0(mesh_3_4_io_in_d_0),
    .io_in_d_1(mesh_3_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_4_io_in_control_1_shift),
    .io_in_id_0(mesh_3_4_io_in_id_0),
    .io_in_id_1(mesh_3_4_io_in_id_1),
    .io_in_last_0(mesh_3_4_io_in_last_0),
    .io_in_last_1(mesh_3_4_io_in_last_1),
    .io_out_a_0(mesh_3_4_io_out_a_0),
    .io_out_a_1(mesh_3_4_io_out_a_1),
    .io_out_c_0(mesh_3_4_io_out_c_0),
    .io_out_c_1(mesh_3_4_io_out_c_1),
    .io_out_b_0(mesh_3_4_io_out_b_0),
    .io_out_b_1(mesh_3_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_4_io_out_control_1_shift),
    .io_out_id_0(mesh_3_4_io_out_id_0),
    .io_out_id_1(mesh_3_4_io_out_id_1),
    .io_out_last_0(mesh_3_4_io_out_last_0),
    .io_out_last_1(mesh_3_4_io_out_last_1),
    .io_in_valid_0(mesh_3_4_io_in_valid_0),
    .io_in_valid_1(mesh_3_4_io_in_valid_1),
    .io_out_valid_0(mesh_3_4_io_out_valid_0),
    .io_out_valid_1(mesh_3_4_io_out_valid_1)
  );
  Tile mesh_3_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_5_clock),
    .io_in_a_0(mesh_3_5_io_in_a_0),
    .io_in_a_1(mesh_3_5_io_in_a_1),
    .io_in_b_0(mesh_3_5_io_in_b_0),
    .io_in_b_1(mesh_3_5_io_in_b_1),
    .io_in_d_0(mesh_3_5_io_in_d_0),
    .io_in_d_1(mesh_3_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_5_io_in_control_1_shift),
    .io_in_id_0(mesh_3_5_io_in_id_0),
    .io_in_id_1(mesh_3_5_io_in_id_1),
    .io_in_last_0(mesh_3_5_io_in_last_0),
    .io_in_last_1(mesh_3_5_io_in_last_1),
    .io_out_a_0(mesh_3_5_io_out_a_0),
    .io_out_a_1(mesh_3_5_io_out_a_1),
    .io_out_c_0(mesh_3_5_io_out_c_0),
    .io_out_c_1(mesh_3_5_io_out_c_1),
    .io_out_b_0(mesh_3_5_io_out_b_0),
    .io_out_b_1(mesh_3_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_5_io_out_control_1_shift),
    .io_out_id_0(mesh_3_5_io_out_id_0),
    .io_out_id_1(mesh_3_5_io_out_id_1),
    .io_out_last_0(mesh_3_5_io_out_last_0),
    .io_out_last_1(mesh_3_5_io_out_last_1),
    .io_in_valid_0(mesh_3_5_io_in_valid_0),
    .io_in_valid_1(mesh_3_5_io_in_valid_1),
    .io_out_valid_0(mesh_3_5_io_out_valid_0),
    .io_out_valid_1(mesh_3_5_io_out_valid_1)
  );
  Tile mesh_3_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_6_clock),
    .io_in_a_0(mesh_3_6_io_in_a_0),
    .io_in_a_1(mesh_3_6_io_in_a_1),
    .io_in_b_0(mesh_3_6_io_in_b_0),
    .io_in_b_1(mesh_3_6_io_in_b_1),
    .io_in_d_0(mesh_3_6_io_in_d_0),
    .io_in_d_1(mesh_3_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_6_io_in_control_1_shift),
    .io_in_id_0(mesh_3_6_io_in_id_0),
    .io_in_id_1(mesh_3_6_io_in_id_1),
    .io_in_last_0(mesh_3_6_io_in_last_0),
    .io_in_last_1(mesh_3_6_io_in_last_1),
    .io_out_a_0(mesh_3_6_io_out_a_0),
    .io_out_a_1(mesh_3_6_io_out_a_1),
    .io_out_c_0(mesh_3_6_io_out_c_0),
    .io_out_c_1(mesh_3_6_io_out_c_1),
    .io_out_b_0(mesh_3_6_io_out_b_0),
    .io_out_b_1(mesh_3_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_6_io_out_control_1_shift),
    .io_out_id_0(mesh_3_6_io_out_id_0),
    .io_out_id_1(mesh_3_6_io_out_id_1),
    .io_out_last_0(mesh_3_6_io_out_last_0),
    .io_out_last_1(mesh_3_6_io_out_last_1),
    .io_in_valid_0(mesh_3_6_io_in_valid_0),
    .io_in_valid_1(mesh_3_6_io_in_valid_1),
    .io_out_valid_0(mesh_3_6_io_out_valid_0),
    .io_out_valid_1(mesh_3_6_io_out_valid_1)
  );
  Tile mesh_3_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_7_clock),
    .io_in_a_0(mesh_3_7_io_in_a_0),
    .io_in_a_1(mesh_3_7_io_in_a_1),
    .io_in_b_0(mesh_3_7_io_in_b_0),
    .io_in_b_1(mesh_3_7_io_in_b_1),
    .io_in_d_0(mesh_3_7_io_in_d_0),
    .io_in_d_1(mesh_3_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_7_io_in_control_1_shift),
    .io_in_id_0(mesh_3_7_io_in_id_0),
    .io_in_id_1(mesh_3_7_io_in_id_1),
    .io_in_last_0(mesh_3_7_io_in_last_0),
    .io_in_last_1(mesh_3_7_io_in_last_1),
    .io_out_a_0(mesh_3_7_io_out_a_0),
    .io_out_a_1(mesh_3_7_io_out_a_1),
    .io_out_c_0(mesh_3_7_io_out_c_0),
    .io_out_c_1(mesh_3_7_io_out_c_1),
    .io_out_b_0(mesh_3_7_io_out_b_0),
    .io_out_b_1(mesh_3_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_7_io_out_control_1_shift),
    .io_out_id_0(mesh_3_7_io_out_id_0),
    .io_out_id_1(mesh_3_7_io_out_id_1),
    .io_out_last_0(mesh_3_7_io_out_last_0),
    .io_out_last_1(mesh_3_7_io_out_last_1),
    .io_in_valid_0(mesh_3_7_io_in_valid_0),
    .io_in_valid_1(mesh_3_7_io_in_valid_1),
    .io_out_valid_0(mesh_3_7_io_out_valid_0),
    .io_out_valid_1(mesh_3_7_io_out_valid_1)
  );
  Tile mesh_3_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_8_clock),
    .io_in_a_0(mesh_3_8_io_in_a_0),
    .io_in_a_1(mesh_3_8_io_in_a_1),
    .io_in_b_0(mesh_3_8_io_in_b_0),
    .io_in_b_1(mesh_3_8_io_in_b_1),
    .io_in_d_0(mesh_3_8_io_in_d_0),
    .io_in_d_1(mesh_3_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_8_io_in_control_1_shift),
    .io_in_id_0(mesh_3_8_io_in_id_0),
    .io_in_id_1(mesh_3_8_io_in_id_1),
    .io_in_last_0(mesh_3_8_io_in_last_0),
    .io_in_last_1(mesh_3_8_io_in_last_1),
    .io_out_a_0(mesh_3_8_io_out_a_0),
    .io_out_a_1(mesh_3_8_io_out_a_1),
    .io_out_c_0(mesh_3_8_io_out_c_0),
    .io_out_c_1(mesh_3_8_io_out_c_1),
    .io_out_b_0(mesh_3_8_io_out_b_0),
    .io_out_b_1(mesh_3_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_8_io_out_control_1_shift),
    .io_out_id_0(mesh_3_8_io_out_id_0),
    .io_out_id_1(mesh_3_8_io_out_id_1),
    .io_out_last_0(mesh_3_8_io_out_last_0),
    .io_out_last_1(mesh_3_8_io_out_last_1),
    .io_in_valid_0(mesh_3_8_io_in_valid_0),
    .io_in_valid_1(mesh_3_8_io_in_valid_1),
    .io_out_valid_0(mesh_3_8_io_out_valid_0),
    .io_out_valid_1(mesh_3_8_io_out_valid_1)
  );
  Tile mesh_3_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_9_clock),
    .io_in_a_0(mesh_3_9_io_in_a_0),
    .io_in_a_1(mesh_3_9_io_in_a_1),
    .io_in_b_0(mesh_3_9_io_in_b_0),
    .io_in_b_1(mesh_3_9_io_in_b_1),
    .io_in_d_0(mesh_3_9_io_in_d_0),
    .io_in_d_1(mesh_3_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_9_io_in_control_1_shift),
    .io_in_id_0(mesh_3_9_io_in_id_0),
    .io_in_id_1(mesh_3_9_io_in_id_1),
    .io_in_last_0(mesh_3_9_io_in_last_0),
    .io_in_last_1(mesh_3_9_io_in_last_1),
    .io_out_a_0(mesh_3_9_io_out_a_0),
    .io_out_a_1(mesh_3_9_io_out_a_1),
    .io_out_c_0(mesh_3_9_io_out_c_0),
    .io_out_c_1(mesh_3_9_io_out_c_1),
    .io_out_b_0(mesh_3_9_io_out_b_0),
    .io_out_b_1(mesh_3_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_9_io_out_control_1_shift),
    .io_out_id_0(mesh_3_9_io_out_id_0),
    .io_out_id_1(mesh_3_9_io_out_id_1),
    .io_out_last_0(mesh_3_9_io_out_last_0),
    .io_out_last_1(mesh_3_9_io_out_last_1),
    .io_in_valid_0(mesh_3_9_io_in_valid_0),
    .io_in_valid_1(mesh_3_9_io_in_valid_1),
    .io_out_valid_0(mesh_3_9_io_out_valid_0),
    .io_out_valid_1(mesh_3_9_io_out_valid_1)
  );
  Tile mesh_3_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_10_clock),
    .io_in_a_0(mesh_3_10_io_in_a_0),
    .io_in_a_1(mesh_3_10_io_in_a_1),
    .io_in_b_0(mesh_3_10_io_in_b_0),
    .io_in_b_1(mesh_3_10_io_in_b_1),
    .io_in_d_0(mesh_3_10_io_in_d_0),
    .io_in_d_1(mesh_3_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_10_io_in_control_1_shift),
    .io_in_id_0(mesh_3_10_io_in_id_0),
    .io_in_id_1(mesh_3_10_io_in_id_1),
    .io_in_last_0(mesh_3_10_io_in_last_0),
    .io_in_last_1(mesh_3_10_io_in_last_1),
    .io_out_a_0(mesh_3_10_io_out_a_0),
    .io_out_a_1(mesh_3_10_io_out_a_1),
    .io_out_c_0(mesh_3_10_io_out_c_0),
    .io_out_c_1(mesh_3_10_io_out_c_1),
    .io_out_b_0(mesh_3_10_io_out_b_0),
    .io_out_b_1(mesh_3_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_10_io_out_control_1_shift),
    .io_out_id_0(mesh_3_10_io_out_id_0),
    .io_out_id_1(mesh_3_10_io_out_id_1),
    .io_out_last_0(mesh_3_10_io_out_last_0),
    .io_out_last_1(mesh_3_10_io_out_last_1),
    .io_in_valid_0(mesh_3_10_io_in_valid_0),
    .io_in_valid_1(mesh_3_10_io_in_valid_1),
    .io_out_valid_0(mesh_3_10_io_out_valid_0),
    .io_out_valid_1(mesh_3_10_io_out_valid_1)
  );
  Tile mesh_3_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_11_clock),
    .io_in_a_0(mesh_3_11_io_in_a_0),
    .io_in_a_1(mesh_3_11_io_in_a_1),
    .io_in_b_0(mesh_3_11_io_in_b_0),
    .io_in_b_1(mesh_3_11_io_in_b_1),
    .io_in_d_0(mesh_3_11_io_in_d_0),
    .io_in_d_1(mesh_3_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_11_io_in_control_1_shift),
    .io_in_id_0(mesh_3_11_io_in_id_0),
    .io_in_id_1(mesh_3_11_io_in_id_1),
    .io_in_last_0(mesh_3_11_io_in_last_0),
    .io_in_last_1(mesh_3_11_io_in_last_1),
    .io_out_a_0(mesh_3_11_io_out_a_0),
    .io_out_a_1(mesh_3_11_io_out_a_1),
    .io_out_c_0(mesh_3_11_io_out_c_0),
    .io_out_c_1(mesh_3_11_io_out_c_1),
    .io_out_b_0(mesh_3_11_io_out_b_0),
    .io_out_b_1(mesh_3_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_11_io_out_control_1_shift),
    .io_out_id_0(mesh_3_11_io_out_id_0),
    .io_out_id_1(mesh_3_11_io_out_id_1),
    .io_out_last_0(mesh_3_11_io_out_last_0),
    .io_out_last_1(mesh_3_11_io_out_last_1),
    .io_in_valid_0(mesh_3_11_io_in_valid_0),
    .io_in_valid_1(mesh_3_11_io_in_valid_1),
    .io_out_valid_0(mesh_3_11_io_out_valid_0),
    .io_out_valid_1(mesh_3_11_io_out_valid_1)
  );
  Tile mesh_3_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_12_clock),
    .io_in_a_0(mesh_3_12_io_in_a_0),
    .io_in_a_1(mesh_3_12_io_in_a_1),
    .io_in_b_0(mesh_3_12_io_in_b_0),
    .io_in_b_1(mesh_3_12_io_in_b_1),
    .io_in_d_0(mesh_3_12_io_in_d_0),
    .io_in_d_1(mesh_3_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_12_io_in_control_1_shift),
    .io_in_id_0(mesh_3_12_io_in_id_0),
    .io_in_id_1(mesh_3_12_io_in_id_1),
    .io_in_last_0(mesh_3_12_io_in_last_0),
    .io_in_last_1(mesh_3_12_io_in_last_1),
    .io_out_a_0(mesh_3_12_io_out_a_0),
    .io_out_a_1(mesh_3_12_io_out_a_1),
    .io_out_c_0(mesh_3_12_io_out_c_0),
    .io_out_c_1(mesh_3_12_io_out_c_1),
    .io_out_b_0(mesh_3_12_io_out_b_0),
    .io_out_b_1(mesh_3_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_12_io_out_control_1_shift),
    .io_out_id_0(mesh_3_12_io_out_id_0),
    .io_out_id_1(mesh_3_12_io_out_id_1),
    .io_out_last_0(mesh_3_12_io_out_last_0),
    .io_out_last_1(mesh_3_12_io_out_last_1),
    .io_in_valid_0(mesh_3_12_io_in_valid_0),
    .io_in_valid_1(mesh_3_12_io_in_valid_1),
    .io_out_valid_0(mesh_3_12_io_out_valid_0),
    .io_out_valid_1(mesh_3_12_io_out_valid_1)
  );
  Tile mesh_3_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_13_clock),
    .io_in_a_0(mesh_3_13_io_in_a_0),
    .io_in_a_1(mesh_3_13_io_in_a_1),
    .io_in_b_0(mesh_3_13_io_in_b_0),
    .io_in_b_1(mesh_3_13_io_in_b_1),
    .io_in_d_0(mesh_3_13_io_in_d_0),
    .io_in_d_1(mesh_3_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_13_io_in_control_1_shift),
    .io_in_id_0(mesh_3_13_io_in_id_0),
    .io_in_id_1(mesh_3_13_io_in_id_1),
    .io_in_last_0(mesh_3_13_io_in_last_0),
    .io_in_last_1(mesh_3_13_io_in_last_1),
    .io_out_a_0(mesh_3_13_io_out_a_0),
    .io_out_a_1(mesh_3_13_io_out_a_1),
    .io_out_c_0(mesh_3_13_io_out_c_0),
    .io_out_c_1(mesh_3_13_io_out_c_1),
    .io_out_b_0(mesh_3_13_io_out_b_0),
    .io_out_b_1(mesh_3_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_13_io_out_control_1_shift),
    .io_out_id_0(mesh_3_13_io_out_id_0),
    .io_out_id_1(mesh_3_13_io_out_id_1),
    .io_out_last_0(mesh_3_13_io_out_last_0),
    .io_out_last_1(mesh_3_13_io_out_last_1),
    .io_in_valid_0(mesh_3_13_io_in_valid_0),
    .io_in_valid_1(mesh_3_13_io_in_valid_1),
    .io_out_valid_0(mesh_3_13_io_out_valid_0),
    .io_out_valid_1(mesh_3_13_io_out_valid_1)
  );
  Tile mesh_3_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_14_clock),
    .io_in_a_0(mesh_3_14_io_in_a_0),
    .io_in_a_1(mesh_3_14_io_in_a_1),
    .io_in_b_0(mesh_3_14_io_in_b_0),
    .io_in_b_1(mesh_3_14_io_in_b_1),
    .io_in_d_0(mesh_3_14_io_in_d_0),
    .io_in_d_1(mesh_3_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_14_io_in_control_1_shift),
    .io_in_id_0(mesh_3_14_io_in_id_0),
    .io_in_id_1(mesh_3_14_io_in_id_1),
    .io_in_last_0(mesh_3_14_io_in_last_0),
    .io_in_last_1(mesh_3_14_io_in_last_1),
    .io_out_a_0(mesh_3_14_io_out_a_0),
    .io_out_a_1(mesh_3_14_io_out_a_1),
    .io_out_c_0(mesh_3_14_io_out_c_0),
    .io_out_c_1(mesh_3_14_io_out_c_1),
    .io_out_b_0(mesh_3_14_io_out_b_0),
    .io_out_b_1(mesh_3_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_14_io_out_control_1_shift),
    .io_out_id_0(mesh_3_14_io_out_id_0),
    .io_out_id_1(mesh_3_14_io_out_id_1),
    .io_out_last_0(mesh_3_14_io_out_last_0),
    .io_out_last_1(mesh_3_14_io_out_last_1),
    .io_in_valid_0(mesh_3_14_io_in_valid_0),
    .io_in_valid_1(mesh_3_14_io_in_valid_1),
    .io_out_valid_0(mesh_3_14_io_out_valid_0),
    .io_out_valid_1(mesh_3_14_io_out_valid_1)
  );
  Tile mesh_3_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_3_15_clock),
    .io_in_a_0(mesh_3_15_io_in_a_0),
    .io_in_a_1(mesh_3_15_io_in_a_1),
    .io_in_b_0(mesh_3_15_io_in_b_0),
    .io_in_b_1(mesh_3_15_io_in_b_1),
    .io_in_d_0(mesh_3_15_io_in_d_0),
    .io_in_d_1(mesh_3_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_3_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_3_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_3_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_3_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_3_15_io_in_control_1_shift),
    .io_in_id_0(mesh_3_15_io_in_id_0),
    .io_in_id_1(mesh_3_15_io_in_id_1),
    .io_in_last_0(mesh_3_15_io_in_last_0),
    .io_in_last_1(mesh_3_15_io_in_last_1),
    .io_out_a_0(mesh_3_15_io_out_a_0),
    .io_out_a_1(mesh_3_15_io_out_a_1),
    .io_out_c_0(mesh_3_15_io_out_c_0),
    .io_out_c_1(mesh_3_15_io_out_c_1),
    .io_out_b_0(mesh_3_15_io_out_b_0),
    .io_out_b_1(mesh_3_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_3_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_3_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_3_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_3_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_3_15_io_out_control_1_shift),
    .io_out_id_0(mesh_3_15_io_out_id_0),
    .io_out_id_1(mesh_3_15_io_out_id_1),
    .io_out_last_0(mesh_3_15_io_out_last_0),
    .io_out_last_1(mesh_3_15_io_out_last_1),
    .io_in_valid_0(mesh_3_15_io_in_valid_0),
    .io_in_valid_1(mesh_3_15_io_in_valid_1),
    .io_out_valid_0(mesh_3_15_io_out_valid_0),
    .io_out_valid_1(mesh_3_15_io_out_valid_1)
  );
  Tile mesh_4_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_0_clock),
    .io_in_a_0(mesh_4_0_io_in_a_0),
    .io_in_a_1(mesh_4_0_io_in_a_1),
    .io_in_b_0(mesh_4_0_io_in_b_0),
    .io_in_b_1(mesh_4_0_io_in_b_1),
    .io_in_d_0(mesh_4_0_io_in_d_0),
    .io_in_d_1(mesh_4_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_0_io_in_control_1_shift),
    .io_in_id_0(mesh_4_0_io_in_id_0),
    .io_in_id_1(mesh_4_0_io_in_id_1),
    .io_in_last_0(mesh_4_0_io_in_last_0),
    .io_in_last_1(mesh_4_0_io_in_last_1),
    .io_out_a_0(mesh_4_0_io_out_a_0),
    .io_out_a_1(mesh_4_0_io_out_a_1),
    .io_out_c_0(mesh_4_0_io_out_c_0),
    .io_out_c_1(mesh_4_0_io_out_c_1),
    .io_out_b_0(mesh_4_0_io_out_b_0),
    .io_out_b_1(mesh_4_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_0_io_out_control_1_shift),
    .io_out_id_0(mesh_4_0_io_out_id_0),
    .io_out_id_1(mesh_4_0_io_out_id_1),
    .io_out_last_0(mesh_4_0_io_out_last_0),
    .io_out_last_1(mesh_4_0_io_out_last_1),
    .io_in_valid_0(mesh_4_0_io_in_valid_0),
    .io_in_valid_1(mesh_4_0_io_in_valid_1),
    .io_out_valid_0(mesh_4_0_io_out_valid_0),
    .io_out_valid_1(mesh_4_0_io_out_valid_1)
  );
  Tile mesh_4_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_1_clock),
    .io_in_a_0(mesh_4_1_io_in_a_0),
    .io_in_a_1(mesh_4_1_io_in_a_1),
    .io_in_b_0(mesh_4_1_io_in_b_0),
    .io_in_b_1(mesh_4_1_io_in_b_1),
    .io_in_d_0(mesh_4_1_io_in_d_0),
    .io_in_d_1(mesh_4_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_1_io_in_control_1_shift),
    .io_in_id_0(mesh_4_1_io_in_id_0),
    .io_in_id_1(mesh_4_1_io_in_id_1),
    .io_in_last_0(mesh_4_1_io_in_last_0),
    .io_in_last_1(mesh_4_1_io_in_last_1),
    .io_out_a_0(mesh_4_1_io_out_a_0),
    .io_out_a_1(mesh_4_1_io_out_a_1),
    .io_out_c_0(mesh_4_1_io_out_c_0),
    .io_out_c_1(mesh_4_1_io_out_c_1),
    .io_out_b_0(mesh_4_1_io_out_b_0),
    .io_out_b_1(mesh_4_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_1_io_out_control_1_shift),
    .io_out_id_0(mesh_4_1_io_out_id_0),
    .io_out_id_1(mesh_4_1_io_out_id_1),
    .io_out_last_0(mesh_4_1_io_out_last_0),
    .io_out_last_1(mesh_4_1_io_out_last_1),
    .io_in_valid_0(mesh_4_1_io_in_valid_0),
    .io_in_valid_1(mesh_4_1_io_in_valid_1),
    .io_out_valid_0(mesh_4_1_io_out_valid_0),
    .io_out_valid_1(mesh_4_1_io_out_valid_1)
  );
  Tile mesh_4_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_2_clock),
    .io_in_a_0(mesh_4_2_io_in_a_0),
    .io_in_a_1(mesh_4_2_io_in_a_1),
    .io_in_b_0(mesh_4_2_io_in_b_0),
    .io_in_b_1(mesh_4_2_io_in_b_1),
    .io_in_d_0(mesh_4_2_io_in_d_0),
    .io_in_d_1(mesh_4_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_2_io_in_control_1_shift),
    .io_in_id_0(mesh_4_2_io_in_id_0),
    .io_in_id_1(mesh_4_2_io_in_id_1),
    .io_in_last_0(mesh_4_2_io_in_last_0),
    .io_in_last_1(mesh_4_2_io_in_last_1),
    .io_out_a_0(mesh_4_2_io_out_a_0),
    .io_out_a_1(mesh_4_2_io_out_a_1),
    .io_out_c_0(mesh_4_2_io_out_c_0),
    .io_out_c_1(mesh_4_2_io_out_c_1),
    .io_out_b_0(mesh_4_2_io_out_b_0),
    .io_out_b_1(mesh_4_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_2_io_out_control_1_shift),
    .io_out_id_0(mesh_4_2_io_out_id_0),
    .io_out_id_1(mesh_4_2_io_out_id_1),
    .io_out_last_0(mesh_4_2_io_out_last_0),
    .io_out_last_1(mesh_4_2_io_out_last_1),
    .io_in_valid_0(mesh_4_2_io_in_valid_0),
    .io_in_valid_1(mesh_4_2_io_in_valid_1),
    .io_out_valid_0(mesh_4_2_io_out_valid_0),
    .io_out_valid_1(mesh_4_2_io_out_valid_1)
  );
  Tile mesh_4_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_3_clock),
    .io_in_a_0(mesh_4_3_io_in_a_0),
    .io_in_a_1(mesh_4_3_io_in_a_1),
    .io_in_b_0(mesh_4_3_io_in_b_0),
    .io_in_b_1(mesh_4_3_io_in_b_1),
    .io_in_d_0(mesh_4_3_io_in_d_0),
    .io_in_d_1(mesh_4_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_3_io_in_control_1_shift),
    .io_in_id_0(mesh_4_3_io_in_id_0),
    .io_in_id_1(mesh_4_3_io_in_id_1),
    .io_in_last_0(mesh_4_3_io_in_last_0),
    .io_in_last_1(mesh_4_3_io_in_last_1),
    .io_out_a_0(mesh_4_3_io_out_a_0),
    .io_out_a_1(mesh_4_3_io_out_a_1),
    .io_out_c_0(mesh_4_3_io_out_c_0),
    .io_out_c_1(mesh_4_3_io_out_c_1),
    .io_out_b_0(mesh_4_3_io_out_b_0),
    .io_out_b_1(mesh_4_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_3_io_out_control_1_shift),
    .io_out_id_0(mesh_4_3_io_out_id_0),
    .io_out_id_1(mesh_4_3_io_out_id_1),
    .io_out_last_0(mesh_4_3_io_out_last_0),
    .io_out_last_1(mesh_4_3_io_out_last_1),
    .io_in_valid_0(mesh_4_3_io_in_valid_0),
    .io_in_valid_1(mesh_4_3_io_in_valid_1),
    .io_out_valid_0(mesh_4_3_io_out_valid_0),
    .io_out_valid_1(mesh_4_3_io_out_valid_1)
  );
  Tile mesh_4_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_4_clock),
    .io_in_a_0(mesh_4_4_io_in_a_0),
    .io_in_a_1(mesh_4_4_io_in_a_1),
    .io_in_b_0(mesh_4_4_io_in_b_0),
    .io_in_b_1(mesh_4_4_io_in_b_1),
    .io_in_d_0(mesh_4_4_io_in_d_0),
    .io_in_d_1(mesh_4_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_4_io_in_control_1_shift),
    .io_in_id_0(mesh_4_4_io_in_id_0),
    .io_in_id_1(mesh_4_4_io_in_id_1),
    .io_in_last_0(mesh_4_4_io_in_last_0),
    .io_in_last_1(mesh_4_4_io_in_last_1),
    .io_out_a_0(mesh_4_4_io_out_a_0),
    .io_out_a_1(mesh_4_4_io_out_a_1),
    .io_out_c_0(mesh_4_4_io_out_c_0),
    .io_out_c_1(mesh_4_4_io_out_c_1),
    .io_out_b_0(mesh_4_4_io_out_b_0),
    .io_out_b_1(mesh_4_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_4_io_out_control_1_shift),
    .io_out_id_0(mesh_4_4_io_out_id_0),
    .io_out_id_1(mesh_4_4_io_out_id_1),
    .io_out_last_0(mesh_4_4_io_out_last_0),
    .io_out_last_1(mesh_4_4_io_out_last_1),
    .io_in_valid_0(mesh_4_4_io_in_valid_0),
    .io_in_valid_1(mesh_4_4_io_in_valid_1),
    .io_out_valid_0(mesh_4_4_io_out_valid_0),
    .io_out_valid_1(mesh_4_4_io_out_valid_1)
  );
  Tile mesh_4_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_5_clock),
    .io_in_a_0(mesh_4_5_io_in_a_0),
    .io_in_a_1(mesh_4_5_io_in_a_1),
    .io_in_b_0(mesh_4_5_io_in_b_0),
    .io_in_b_1(mesh_4_5_io_in_b_1),
    .io_in_d_0(mesh_4_5_io_in_d_0),
    .io_in_d_1(mesh_4_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_5_io_in_control_1_shift),
    .io_in_id_0(mesh_4_5_io_in_id_0),
    .io_in_id_1(mesh_4_5_io_in_id_1),
    .io_in_last_0(mesh_4_5_io_in_last_0),
    .io_in_last_1(mesh_4_5_io_in_last_1),
    .io_out_a_0(mesh_4_5_io_out_a_0),
    .io_out_a_1(mesh_4_5_io_out_a_1),
    .io_out_c_0(mesh_4_5_io_out_c_0),
    .io_out_c_1(mesh_4_5_io_out_c_1),
    .io_out_b_0(mesh_4_5_io_out_b_0),
    .io_out_b_1(mesh_4_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_5_io_out_control_1_shift),
    .io_out_id_0(mesh_4_5_io_out_id_0),
    .io_out_id_1(mesh_4_5_io_out_id_1),
    .io_out_last_0(mesh_4_5_io_out_last_0),
    .io_out_last_1(mesh_4_5_io_out_last_1),
    .io_in_valid_0(mesh_4_5_io_in_valid_0),
    .io_in_valid_1(mesh_4_5_io_in_valid_1),
    .io_out_valid_0(mesh_4_5_io_out_valid_0),
    .io_out_valid_1(mesh_4_5_io_out_valid_1)
  );
  Tile mesh_4_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_6_clock),
    .io_in_a_0(mesh_4_6_io_in_a_0),
    .io_in_a_1(mesh_4_6_io_in_a_1),
    .io_in_b_0(mesh_4_6_io_in_b_0),
    .io_in_b_1(mesh_4_6_io_in_b_1),
    .io_in_d_0(mesh_4_6_io_in_d_0),
    .io_in_d_1(mesh_4_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_6_io_in_control_1_shift),
    .io_in_id_0(mesh_4_6_io_in_id_0),
    .io_in_id_1(mesh_4_6_io_in_id_1),
    .io_in_last_0(mesh_4_6_io_in_last_0),
    .io_in_last_1(mesh_4_6_io_in_last_1),
    .io_out_a_0(mesh_4_6_io_out_a_0),
    .io_out_a_1(mesh_4_6_io_out_a_1),
    .io_out_c_0(mesh_4_6_io_out_c_0),
    .io_out_c_1(mesh_4_6_io_out_c_1),
    .io_out_b_0(mesh_4_6_io_out_b_0),
    .io_out_b_1(mesh_4_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_6_io_out_control_1_shift),
    .io_out_id_0(mesh_4_6_io_out_id_0),
    .io_out_id_1(mesh_4_6_io_out_id_1),
    .io_out_last_0(mesh_4_6_io_out_last_0),
    .io_out_last_1(mesh_4_6_io_out_last_1),
    .io_in_valid_0(mesh_4_6_io_in_valid_0),
    .io_in_valid_1(mesh_4_6_io_in_valid_1),
    .io_out_valid_0(mesh_4_6_io_out_valid_0),
    .io_out_valid_1(mesh_4_6_io_out_valid_1)
  );
  Tile mesh_4_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_7_clock),
    .io_in_a_0(mesh_4_7_io_in_a_0),
    .io_in_a_1(mesh_4_7_io_in_a_1),
    .io_in_b_0(mesh_4_7_io_in_b_0),
    .io_in_b_1(mesh_4_7_io_in_b_1),
    .io_in_d_0(mesh_4_7_io_in_d_0),
    .io_in_d_1(mesh_4_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_7_io_in_control_1_shift),
    .io_in_id_0(mesh_4_7_io_in_id_0),
    .io_in_id_1(mesh_4_7_io_in_id_1),
    .io_in_last_0(mesh_4_7_io_in_last_0),
    .io_in_last_1(mesh_4_7_io_in_last_1),
    .io_out_a_0(mesh_4_7_io_out_a_0),
    .io_out_a_1(mesh_4_7_io_out_a_1),
    .io_out_c_0(mesh_4_7_io_out_c_0),
    .io_out_c_1(mesh_4_7_io_out_c_1),
    .io_out_b_0(mesh_4_7_io_out_b_0),
    .io_out_b_1(mesh_4_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_7_io_out_control_1_shift),
    .io_out_id_0(mesh_4_7_io_out_id_0),
    .io_out_id_1(mesh_4_7_io_out_id_1),
    .io_out_last_0(mesh_4_7_io_out_last_0),
    .io_out_last_1(mesh_4_7_io_out_last_1),
    .io_in_valid_0(mesh_4_7_io_in_valid_0),
    .io_in_valid_1(mesh_4_7_io_in_valid_1),
    .io_out_valid_0(mesh_4_7_io_out_valid_0),
    .io_out_valid_1(mesh_4_7_io_out_valid_1)
  );
  Tile mesh_4_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_8_clock),
    .io_in_a_0(mesh_4_8_io_in_a_0),
    .io_in_a_1(mesh_4_8_io_in_a_1),
    .io_in_b_0(mesh_4_8_io_in_b_0),
    .io_in_b_1(mesh_4_8_io_in_b_1),
    .io_in_d_0(mesh_4_8_io_in_d_0),
    .io_in_d_1(mesh_4_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_8_io_in_control_1_shift),
    .io_in_id_0(mesh_4_8_io_in_id_0),
    .io_in_id_1(mesh_4_8_io_in_id_1),
    .io_in_last_0(mesh_4_8_io_in_last_0),
    .io_in_last_1(mesh_4_8_io_in_last_1),
    .io_out_a_0(mesh_4_8_io_out_a_0),
    .io_out_a_1(mesh_4_8_io_out_a_1),
    .io_out_c_0(mesh_4_8_io_out_c_0),
    .io_out_c_1(mesh_4_8_io_out_c_1),
    .io_out_b_0(mesh_4_8_io_out_b_0),
    .io_out_b_1(mesh_4_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_8_io_out_control_1_shift),
    .io_out_id_0(mesh_4_8_io_out_id_0),
    .io_out_id_1(mesh_4_8_io_out_id_1),
    .io_out_last_0(mesh_4_8_io_out_last_0),
    .io_out_last_1(mesh_4_8_io_out_last_1),
    .io_in_valid_0(mesh_4_8_io_in_valid_0),
    .io_in_valid_1(mesh_4_8_io_in_valid_1),
    .io_out_valid_0(mesh_4_8_io_out_valid_0),
    .io_out_valid_1(mesh_4_8_io_out_valid_1)
  );
  Tile mesh_4_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_9_clock),
    .io_in_a_0(mesh_4_9_io_in_a_0),
    .io_in_a_1(mesh_4_9_io_in_a_1),
    .io_in_b_0(mesh_4_9_io_in_b_0),
    .io_in_b_1(mesh_4_9_io_in_b_1),
    .io_in_d_0(mesh_4_9_io_in_d_0),
    .io_in_d_1(mesh_4_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_9_io_in_control_1_shift),
    .io_in_id_0(mesh_4_9_io_in_id_0),
    .io_in_id_1(mesh_4_9_io_in_id_1),
    .io_in_last_0(mesh_4_9_io_in_last_0),
    .io_in_last_1(mesh_4_9_io_in_last_1),
    .io_out_a_0(mesh_4_9_io_out_a_0),
    .io_out_a_1(mesh_4_9_io_out_a_1),
    .io_out_c_0(mesh_4_9_io_out_c_0),
    .io_out_c_1(mesh_4_9_io_out_c_1),
    .io_out_b_0(mesh_4_9_io_out_b_0),
    .io_out_b_1(mesh_4_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_9_io_out_control_1_shift),
    .io_out_id_0(mesh_4_9_io_out_id_0),
    .io_out_id_1(mesh_4_9_io_out_id_1),
    .io_out_last_0(mesh_4_9_io_out_last_0),
    .io_out_last_1(mesh_4_9_io_out_last_1),
    .io_in_valid_0(mesh_4_9_io_in_valid_0),
    .io_in_valid_1(mesh_4_9_io_in_valid_1),
    .io_out_valid_0(mesh_4_9_io_out_valid_0),
    .io_out_valid_1(mesh_4_9_io_out_valid_1)
  );
  Tile mesh_4_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_10_clock),
    .io_in_a_0(mesh_4_10_io_in_a_0),
    .io_in_a_1(mesh_4_10_io_in_a_1),
    .io_in_b_0(mesh_4_10_io_in_b_0),
    .io_in_b_1(mesh_4_10_io_in_b_1),
    .io_in_d_0(mesh_4_10_io_in_d_0),
    .io_in_d_1(mesh_4_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_10_io_in_control_1_shift),
    .io_in_id_0(mesh_4_10_io_in_id_0),
    .io_in_id_1(mesh_4_10_io_in_id_1),
    .io_in_last_0(mesh_4_10_io_in_last_0),
    .io_in_last_1(mesh_4_10_io_in_last_1),
    .io_out_a_0(mesh_4_10_io_out_a_0),
    .io_out_a_1(mesh_4_10_io_out_a_1),
    .io_out_c_0(mesh_4_10_io_out_c_0),
    .io_out_c_1(mesh_4_10_io_out_c_1),
    .io_out_b_0(mesh_4_10_io_out_b_0),
    .io_out_b_1(mesh_4_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_10_io_out_control_1_shift),
    .io_out_id_0(mesh_4_10_io_out_id_0),
    .io_out_id_1(mesh_4_10_io_out_id_1),
    .io_out_last_0(mesh_4_10_io_out_last_0),
    .io_out_last_1(mesh_4_10_io_out_last_1),
    .io_in_valid_0(mesh_4_10_io_in_valid_0),
    .io_in_valid_1(mesh_4_10_io_in_valid_1),
    .io_out_valid_0(mesh_4_10_io_out_valid_0),
    .io_out_valid_1(mesh_4_10_io_out_valid_1)
  );
  Tile mesh_4_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_11_clock),
    .io_in_a_0(mesh_4_11_io_in_a_0),
    .io_in_a_1(mesh_4_11_io_in_a_1),
    .io_in_b_0(mesh_4_11_io_in_b_0),
    .io_in_b_1(mesh_4_11_io_in_b_1),
    .io_in_d_0(mesh_4_11_io_in_d_0),
    .io_in_d_1(mesh_4_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_11_io_in_control_1_shift),
    .io_in_id_0(mesh_4_11_io_in_id_0),
    .io_in_id_1(mesh_4_11_io_in_id_1),
    .io_in_last_0(mesh_4_11_io_in_last_0),
    .io_in_last_1(mesh_4_11_io_in_last_1),
    .io_out_a_0(mesh_4_11_io_out_a_0),
    .io_out_a_1(mesh_4_11_io_out_a_1),
    .io_out_c_0(mesh_4_11_io_out_c_0),
    .io_out_c_1(mesh_4_11_io_out_c_1),
    .io_out_b_0(mesh_4_11_io_out_b_0),
    .io_out_b_1(mesh_4_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_11_io_out_control_1_shift),
    .io_out_id_0(mesh_4_11_io_out_id_0),
    .io_out_id_1(mesh_4_11_io_out_id_1),
    .io_out_last_0(mesh_4_11_io_out_last_0),
    .io_out_last_1(mesh_4_11_io_out_last_1),
    .io_in_valid_0(mesh_4_11_io_in_valid_0),
    .io_in_valid_1(mesh_4_11_io_in_valid_1),
    .io_out_valid_0(mesh_4_11_io_out_valid_0),
    .io_out_valid_1(mesh_4_11_io_out_valid_1)
  );
  Tile mesh_4_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_12_clock),
    .io_in_a_0(mesh_4_12_io_in_a_0),
    .io_in_a_1(mesh_4_12_io_in_a_1),
    .io_in_b_0(mesh_4_12_io_in_b_0),
    .io_in_b_1(mesh_4_12_io_in_b_1),
    .io_in_d_0(mesh_4_12_io_in_d_0),
    .io_in_d_1(mesh_4_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_12_io_in_control_1_shift),
    .io_in_id_0(mesh_4_12_io_in_id_0),
    .io_in_id_1(mesh_4_12_io_in_id_1),
    .io_in_last_0(mesh_4_12_io_in_last_0),
    .io_in_last_1(mesh_4_12_io_in_last_1),
    .io_out_a_0(mesh_4_12_io_out_a_0),
    .io_out_a_1(mesh_4_12_io_out_a_1),
    .io_out_c_0(mesh_4_12_io_out_c_0),
    .io_out_c_1(mesh_4_12_io_out_c_1),
    .io_out_b_0(mesh_4_12_io_out_b_0),
    .io_out_b_1(mesh_4_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_12_io_out_control_1_shift),
    .io_out_id_0(mesh_4_12_io_out_id_0),
    .io_out_id_1(mesh_4_12_io_out_id_1),
    .io_out_last_0(mesh_4_12_io_out_last_0),
    .io_out_last_1(mesh_4_12_io_out_last_1),
    .io_in_valid_0(mesh_4_12_io_in_valid_0),
    .io_in_valid_1(mesh_4_12_io_in_valid_1),
    .io_out_valid_0(mesh_4_12_io_out_valid_0),
    .io_out_valid_1(mesh_4_12_io_out_valid_1)
  );
  Tile mesh_4_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_13_clock),
    .io_in_a_0(mesh_4_13_io_in_a_0),
    .io_in_a_1(mesh_4_13_io_in_a_1),
    .io_in_b_0(mesh_4_13_io_in_b_0),
    .io_in_b_1(mesh_4_13_io_in_b_1),
    .io_in_d_0(mesh_4_13_io_in_d_0),
    .io_in_d_1(mesh_4_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_13_io_in_control_1_shift),
    .io_in_id_0(mesh_4_13_io_in_id_0),
    .io_in_id_1(mesh_4_13_io_in_id_1),
    .io_in_last_0(mesh_4_13_io_in_last_0),
    .io_in_last_1(mesh_4_13_io_in_last_1),
    .io_out_a_0(mesh_4_13_io_out_a_0),
    .io_out_a_1(mesh_4_13_io_out_a_1),
    .io_out_c_0(mesh_4_13_io_out_c_0),
    .io_out_c_1(mesh_4_13_io_out_c_1),
    .io_out_b_0(mesh_4_13_io_out_b_0),
    .io_out_b_1(mesh_4_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_13_io_out_control_1_shift),
    .io_out_id_0(mesh_4_13_io_out_id_0),
    .io_out_id_1(mesh_4_13_io_out_id_1),
    .io_out_last_0(mesh_4_13_io_out_last_0),
    .io_out_last_1(mesh_4_13_io_out_last_1),
    .io_in_valid_0(mesh_4_13_io_in_valid_0),
    .io_in_valid_1(mesh_4_13_io_in_valid_1),
    .io_out_valid_0(mesh_4_13_io_out_valid_0),
    .io_out_valid_1(mesh_4_13_io_out_valid_1)
  );
  Tile mesh_4_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_14_clock),
    .io_in_a_0(mesh_4_14_io_in_a_0),
    .io_in_a_1(mesh_4_14_io_in_a_1),
    .io_in_b_0(mesh_4_14_io_in_b_0),
    .io_in_b_1(mesh_4_14_io_in_b_1),
    .io_in_d_0(mesh_4_14_io_in_d_0),
    .io_in_d_1(mesh_4_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_14_io_in_control_1_shift),
    .io_in_id_0(mesh_4_14_io_in_id_0),
    .io_in_id_1(mesh_4_14_io_in_id_1),
    .io_in_last_0(mesh_4_14_io_in_last_0),
    .io_in_last_1(mesh_4_14_io_in_last_1),
    .io_out_a_0(mesh_4_14_io_out_a_0),
    .io_out_a_1(mesh_4_14_io_out_a_1),
    .io_out_c_0(mesh_4_14_io_out_c_0),
    .io_out_c_1(mesh_4_14_io_out_c_1),
    .io_out_b_0(mesh_4_14_io_out_b_0),
    .io_out_b_1(mesh_4_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_14_io_out_control_1_shift),
    .io_out_id_0(mesh_4_14_io_out_id_0),
    .io_out_id_1(mesh_4_14_io_out_id_1),
    .io_out_last_0(mesh_4_14_io_out_last_0),
    .io_out_last_1(mesh_4_14_io_out_last_1),
    .io_in_valid_0(mesh_4_14_io_in_valid_0),
    .io_in_valid_1(mesh_4_14_io_in_valid_1),
    .io_out_valid_0(mesh_4_14_io_out_valid_0),
    .io_out_valid_1(mesh_4_14_io_out_valid_1)
  );
  Tile mesh_4_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_4_15_clock),
    .io_in_a_0(mesh_4_15_io_in_a_0),
    .io_in_a_1(mesh_4_15_io_in_a_1),
    .io_in_b_0(mesh_4_15_io_in_b_0),
    .io_in_b_1(mesh_4_15_io_in_b_1),
    .io_in_d_0(mesh_4_15_io_in_d_0),
    .io_in_d_1(mesh_4_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_4_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_4_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_4_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_4_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_4_15_io_in_control_1_shift),
    .io_in_id_0(mesh_4_15_io_in_id_0),
    .io_in_id_1(mesh_4_15_io_in_id_1),
    .io_in_last_0(mesh_4_15_io_in_last_0),
    .io_in_last_1(mesh_4_15_io_in_last_1),
    .io_out_a_0(mesh_4_15_io_out_a_0),
    .io_out_a_1(mesh_4_15_io_out_a_1),
    .io_out_c_0(mesh_4_15_io_out_c_0),
    .io_out_c_1(mesh_4_15_io_out_c_1),
    .io_out_b_0(mesh_4_15_io_out_b_0),
    .io_out_b_1(mesh_4_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_4_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_4_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_4_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_4_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_4_15_io_out_control_1_shift),
    .io_out_id_0(mesh_4_15_io_out_id_0),
    .io_out_id_1(mesh_4_15_io_out_id_1),
    .io_out_last_0(mesh_4_15_io_out_last_0),
    .io_out_last_1(mesh_4_15_io_out_last_1),
    .io_in_valid_0(mesh_4_15_io_in_valid_0),
    .io_in_valid_1(mesh_4_15_io_in_valid_1),
    .io_out_valid_0(mesh_4_15_io_out_valid_0),
    .io_out_valid_1(mesh_4_15_io_out_valid_1)
  );
  Tile mesh_5_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_0_clock),
    .io_in_a_0(mesh_5_0_io_in_a_0),
    .io_in_a_1(mesh_5_0_io_in_a_1),
    .io_in_b_0(mesh_5_0_io_in_b_0),
    .io_in_b_1(mesh_5_0_io_in_b_1),
    .io_in_d_0(mesh_5_0_io_in_d_0),
    .io_in_d_1(mesh_5_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_0_io_in_control_1_shift),
    .io_in_id_0(mesh_5_0_io_in_id_0),
    .io_in_id_1(mesh_5_0_io_in_id_1),
    .io_in_last_0(mesh_5_0_io_in_last_0),
    .io_in_last_1(mesh_5_0_io_in_last_1),
    .io_out_a_0(mesh_5_0_io_out_a_0),
    .io_out_a_1(mesh_5_0_io_out_a_1),
    .io_out_c_0(mesh_5_0_io_out_c_0),
    .io_out_c_1(mesh_5_0_io_out_c_1),
    .io_out_b_0(mesh_5_0_io_out_b_0),
    .io_out_b_1(mesh_5_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_0_io_out_control_1_shift),
    .io_out_id_0(mesh_5_0_io_out_id_0),
    .io_out_id_1(mesh_5_0_io_out_id_1),
    .io_out_last_0(mesh_5_0_io_out_last_0),
    .io_out_last_1(mesh_5_0_io_out_last_1),
    .io_in_valid_0(mesh_5_0_io_in_valid_0),
    .io_in_valid_1(mesh_5_0_io_in_valid_1),
    .io_out_valid_0(mesh_5_0_io_out_valid_0),
    .io_out_valid_1(mesh_5_0_io_out_valid_1)
  );
  Tile mesh_5_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_1_clock),
    .io_in_a_0(mesh_5_1_io_in_a_0),
    .io_in_a_1(mesh_5_1_io_in_a_1),
    .io_in_b_0(mesh_5_1_io_in_b_0),
    .io_in_b_1(mesh_5_1_io_in_b_1),
    .io_in_d_0(mesh_5_1_io_in_d_0),
    .io_in_d_1(mesh_5_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_1_io_in_control_1_shift),
    .io_in_id_0(mesh_5_1_io_in_id_0),
    .io_in_id_1(mesh_5_1_io_in_id_1),
    .io_in_last_0(mesh_5_1_io_in_last_0),
    .io_in_last_1(mesh_5_1_io_in_last_1),
    .io_out_a_0(mesh_5_1_io_out_a_0),
    .io_out_a_1(mesh_5_1_io_out_a_1),
    .io_out_c_0(mesh_5_1_io_out_c_0),
    .io_out_c_1(mesh_5_1_io_out_c_1),
    .io_out_b_0(mesh_5_1_io_out_b_0),
    .io_out_b_1(mesh_5_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_1_io_out_control_1_shift),
    .io_out_id_0(mesh_5_1_io_out_id_0),
    .io_out_id_1(mesh_5_1_io_out_id_1),
    .io_out_last_0(mesh_5_1_io_out_last_0),
    .io_out_last_1(mesh_5_1_io_out_last_1),
    .io_in_valid_0(mesh_5_1_io_in_valid_0),
    .io_in_valid_1(mesh_5_1_io_in_valid_1),
    .io_out_valid_0(mesh_5_1_io_out_valid_0),
    .io_out_valid_1(mesh_5_1_io_out_valid_1)
  );
  Tile mesh_5_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_2_clock),
    .io_in_a_0(mesh_5_2_io_in_a_0),
    .io_in_a_1(mesh_5_2_io_in_a_1),
    .io_in_b_0(mesh_5_2_io_in_b_0),
    .io_in_b_1(mesh_5_2_io_in_b_1),
    .io_in_d_0(mesh_5_2_io_in_d_0),
    .io_in_d_1(mesh_5_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_2_io_in_control_1_shift),
    .io_in_id_0(mesh_5_2_io_in_id_0),
    .io_in_id_1(mesh_5_2_io_in_id_1),
    .io_in_last_0(mesh_5_2_io_in_last_0),
    .io_in_last_1(mesh_5_2_io_in_last_1),
    .io_out_a_0(mesh_5_2_io_out_a_0),
    .io_out_a_1(mesh_5_2_io_out_a_1),
    .io_out_c_0(mesh_5_2_io_out_c_0),
    .io_out_c_1(mesh_5_2_io_out_c_1),
    .io_out_b_0(mesh_5_2_io_out_b_0),
    .io_out_b_1(mesh_5_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_2_io_out_control_1_shift),
    .io_out_id_0(mesh_5_2_io_out_id_0),
    .io_out_id_1(mesh_5_2_io_out_id_1),
    .io_out_last_0(mesh_5_2_io_out_last_0),
    .io_out_last_1(mesh_5_2_io_out_last_1),
    .io_in_valid_0(mesh_5_2_io_in_valid_0),
    .io_in_valid_1(mesh_5_2_io_in_valid_1),
    .io_out_valid_0(mesh_5_2_io_out_valid_0),
    .io_out_valid_1(mesh_5_2_io_out_valid_1)
  );
  Tile mesh_5_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_3_clock),
    .io_in_a_0(mesh_5_3_io_in_a_0),
    .io_in_a_1(mesh_5_3_io_in_a_1),
    .io_in_b_0(mesh_5_3_io_in_b_0),
    .io_in_b_1(mesh_5_3_io_in_b_1),
    .io_in_d_0(mesh_5_3_io_in_d_0),
    .io_in_d_1(mesh_5_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_3_io_in_control_1_shift),
    .io_in_id_0(mesh_5_3_io_in_id_0),
    .io_in_id_1(mesh_5_3_io_in_id_1),
    .io_in_last_0(mesh_5_3_io_in_last_0),
    .io_in_last_1(mesh_5_3_io_in_last_1),
    .io_out_a_0(mesh_5_3_io_out_a_0),
    .io_out_a_1(mesh_5_3_io_out_a_1),
    .io_out_c_0(mesh_5_3_io_out_c_0),
    .io_out_c_1(mesh_5_3_io_out_c_1),
    .io_out_b_0(mesh_5_3_io_out_b_0),
    .io_out_b_1(mesh_5_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_3_io_out_control_1_shift),
    .io_out_id_0(mesh_5_3_io_out_id_0),
    .io_out_id_1(mesh_5_3_io_out_id_1),
    .io_out_last_0(mesh_5_3_io_out_last_0),
    .io_out_last_1(mesh_5_3_io_out_last_1),
    .io_in_valid_0(mesh_5_3_io_in_valid_0),
    .io_in_valid_1(mesh_5_3_io_in_valid_1),
    .io_out_valid_0(mesh_5_3_io_out_valid_0),
    .io_out_valid_1(mesh_5_3_io_out_valid_1)
  );
  Tile mesh_5_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_4_clock),
    .io_in_a_0(mesh_5_4_io_in_a_0),
    .io_in_a_1(mesh_5_4_io_in_a_1),
    .io_in_b_0(mesh_5_4_io_in_b_0),
    .io_in_b_1(mesh_5_4_io_in_b_1),
    .io_in_d_0(mesh_5_4_io_in_d_0),
    .io_in_d_1(mesh_5_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_4_io_in_control_1_shift),
    .io_in_id_0(mesh_5_4_io_in_id_0),
    .io_in_id_1(mesh_5_4_io_in_id_1),
    .io_in_last_0(mesh_5_4_io_in_last_0),
    .io_in_last_1(mesh_5_4_io_in_last_1),
    .io_out_a_0(mesh_5_4_io_out_a_0),
    .io_out_a_1(mesh_5_4_io_out_a_1),
    .io_out_c_0(mesh_5_4_io_out_c_0),
    .io_out_c_1(mesh_5_4_io_out_c_1),
    .io_out_b_0(mesh_5_4_io_out_b_0),
    .io_out_b_1(mesh_5_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_4_io_out_control_1_shift),
    .io_out_id_0(mesh_5_4_io_out_id_0),
    .io_out_id_1(mesh_5_4_io_out_id_1),
    .io_out_last_0(mesh_5_4_io_out_last_0),
    .io_out_last_1(mesh_5_4_io_out_last_1),
    .io_in_valid_0(mesh_5_4_io_in_valid_0),
    .io_in_valid_1(mesh_5_4_io_in_valid_1),
    .io_out_valid_0(mesh_5_4_io_out_valid_0),
    .io_out_valid_1(mesh_5_4_io_out_valid_1)
  );
  Tile mesh_5_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_5_clock),
    .io_in_a_0(mesh_5_5_io_in_a_0),
    .io_in_a_1(mesh_5_5_io_in_a_1),
    .io_in_b_0(mesh_5_5_io_in_b_0),
    .io_in_b_1(mesh_5_5_io_in_b_1),
    .io_in_d_0(mesh_5_5_io_in_d_0),
    .io_in_d_1(mesh_5_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_5_io_in_control_1_shift),
    .io_in_id_0(mesh_5_5_io_in_id_0),
    .io_in_id_1(mesh_5_5_io_in_id_1),
    .io_in_last_0(mesh_5_5_io_in_last_0),
    .io_in_last_1(mesh_5_5_io_in_last_1),
    .io_out_a_0(mesh_5_5_io_out_a_0),
    .io_out_a_1(mesh_5_5_io_out_a_1),
    .io_out_c_0(mesh_5_5_io_out_c_0),
    .io_out_c_1(mesh_5_5_io_out_c_1),
    .io_out_b_0(mesh_5_5_io_out_b_0),
    .io_out_b_1(mesh_5_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_5_io_out_control_1_shift),
    .io_out_id_0(mesh_5_5_io_out_id_0),
    .io_out_id_1(mesh_5_5_io_out_id_1),
    .io_out_last_0(mesh_5_5_io_out_last_0),
    .io_out_last_1(mesh_5_5_io_out_last_1),
    .io_in_valid_0(mesh_5_5_io_in_valid_0),
    .io_in_valid_1(mesh_5_5_io_in_valid_1),
    .io_out_valid_0(mesh_5_5_io_out_valid_0),
    .io_out_valid_1(mesh_5_5_io_out_valid_1)
  );
  Tile mesh_5_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_6_clock),
    .io_in_a_0(mesh_5_6_io_in_a_0),
    .io_in_a_1(mesh_5_6_io_in_a_1),
    .io_in_b_0(mesh_5_6_io_in_b_0),
    .io_in_b_1(mesh_5_6_io_in_b_1),
    .io_in_d_0(mesh_5_6_io_in_d_0),
    .io_in_d_1(mesh_5_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_6_io_in_control_1_shift),
    .io_in_id_0(mesh_5_6_io_in_id_0),
    .io_in_id_1(mesh_5_6_io_in_id_1),
    .io_in_last_0(mesh_5_6_io_in_last_0),
    .io_in_last_1(mesh_5_6_io_in_last_1),
    .io_out_a_0(mesh_5_6_io_out_a_0),
    .io_out_a_1(mesh_5_6_io_out_a_1),
    .io_out_c_0(mesh_5_6_io_out_c_0),
    .io_out_c_1(mesh_5_6_io_out_c_1),
    .io_out_b_0(mesh_5_6_io_out_b_0),
    .io_out_b_1(mesh_5_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_6_io_out_control_1_shift),
    .io_out_id_0(mesh_5_6_io_out_id_0),
    .io_out_id_1(mesh_5_6_io_out_id_1),
    .io_out_last_0(mesh_5_6_io_out_last_0),
    .io_out_last_1(mesh_5_6_io_out_last_1),
    .io_in_valid_0(mesh_5_6_io_in_valid_0),
    .io_in_valid_1(mesh_5_6_io_in_valid_1),
    .io_out_valid_0(mesh_5_6_io_out_valid_0),
    .io_out_valid_1(mesh_5_6_io_out_valid_1)
  );
  Tile mesh_5_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_7_clock),
    .io_in_a_0(mesh_5_7_io_in_a_0),
    .io_in_a_1(mesh_5_7_io_in_a_1),
    .io_in_b_0(mesh_5_7_io_in_b_0),
    .io_in_b_1(mesh_5_7_io_in_b_1),
    .io_in_d_0(mesh_5_7_io_in_d_0),
    .io_in_d_1(mesh_5_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_7_io_in_control_1_shift),
    .io_in_id_0(mesh_5_7_io_in_id_0),
    .io_in_id_1(mesh_5_7_io_in_id_1),
    .io_in_last_0(mesh_5_7_io_in_last_0),
    .io_in_last_1(mesh_5_7_io_in_last_1),
    .io_out_a_0(mesh_5_7_io_out_a_0),
    .io_out_a_1(mesh_5_7_io_out_a_1),
    .io_out_c_0(mesh_5_7_io_out_c_0),
    .io_out_c_1(mesh_5_7_io_out_c_1),
    .io_out_b_0(mesh_5_7_io_out_b_0),
    .io_out_b_1(mesh_5_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_7_io_out_control_1_shift),
    .io_out_id_0(mesh_5_7_io_out_id_0),
    .io_out_id_1(mesh_5_7_io_out_id_1),
    .io_out_last_0(mesh_5_7_io_out_last_0),
    .io_out_last_1(mesh_5_7_io_out_last_1),
    .io_in_valid_0(mesh_5_7_io_in_valid_0),
    .io_in_valid_1(mesh_5_7_io_in_valid_1),
    .io_out_valid_0(mesh_5_7_io_out_valid_0),
    .io_out_valid_1(mesh_5_7_io_out_valid_1)
  );
  Tile mesh_5_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_8_clock),
    .io_in_a_0(mesh_5_8_io_in_a_0),
    .io_in_a_1(mesh_5_8_io_in_a_1),
    .io_in_b_0(mesh_5_8_io_in_b_0),
    .io_in_b_1(mesh_5_8_io_in_b_1),
    .io_in_d_0(mesh_5_8_io_in_d_0),
    .io_in_d_1(mesh_5_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_8_io_in_control_1_shift),
    .io_in_id_0(mesh_5_8_io_in_id_0),
    .io_in_id_1(mesh_5_8_io_in_id_1),
    .io_in_last_0(mesh_5_8_io_in_last_0),
    .io_in_last_1(mesh_5_8_io_in_last_1),
    .io_out_a_0(mesh_5_8_io_out_a_0),
    .io_out_a_1(mesh_5_8_io_out_a_1),
    .io_out_c_0(mesh_5_8_io_out_c_0),
    .io_out_c_1(mesh_5_8_io_out_c_1),
    .io_out_b_0(mesh_5_8_io_out_b_0),
    .io_out_b_1(mesh_5_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_8_io_out_control_1_shift),
    .io_out_id_0(mesh_5_8_io_out_id_0),
    .io_out_id_1(mesh_5_8_io_out_id_1),
    .io_out_last_0(mesh_5_8_io_out_last_0),
    .io_out_last_1(mesh_5_8_io_out_last_1),
    .io_in_valid_0(mesh_5_8_io_in_valid_0),
    .io_in_valid_1(mesh_5_8_io_in_valid_1),
    .io_out_valid_0(mesh_5_8_io_out_valid_0),
    .io_out_valid_1(mesh_5_8_io_out_valid_1)
  );
  Tile mesh_5_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_9_clock),
    .io_in_a_0(mesh_5_9_io_in_a_0),
    .io_in_a_1(mesh_5_9_io_in_a_1),
    .io_in_b_0(mesh_5_9_io_in_b_0),
    .io_in_b_1(mesh_5_9_io_in_b_1),
    .io_in_d_0(mesh_5_9_io_in_d_0),
    .io_in_d_1(mesh_5_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_9_io_in_control_1_shift),
    .io_in_id_0(mesh_5_9_io_in_id_0),
    .io_in_id_1(mesh_5_9_io_in_id_1),
    .io_in_last_0(mesh_5_9_io_in_last_0),
    .io_in_last_1(mesh_5_9_io_in_last_1),
    .io_out_a_0(mesh_5_9_io_out_a_0),
    .io_out_a_1(mesh_5_9_io_out_a_1),
    .io_out_c_0(mesh_5_9_io_out_c_0),
    .io_out_c_1(mesh_5_9_io_out_c_1),
    .io_out_b_0(mesh_5_9_io_out_b_0),
    .io_out_b_1(mesh_5_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_9_io_out_control_1_shift),
    .io_out_id_0(mesh_5_9_io_out_id_0),
    .io_out_id_1(mesh_5_9_io_out_id_1),
    .io_out_last_0(mesh_5_9_io_out_last_0),
    .io_out_last_1(mesh_5_9_io_out_last_1),
    .io_in_valid_0(mesh_5_9_io_in_valid_0),
    .io_in_valid_1(mesh_5_9_io_in_valid_1),
    .io_out_valid_0(mesh_5_9_io_out_valid_0),
    .io_out_valid_1(mesh_5_9_io_out_valid_1)
  );
  Tile mesh_5_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_10_clock),
    .io_in_a_0(mesh_5_10_io_in_a_0),
    .io_in_a_1(mesh_5_10_io_in_a_1),
    .io_in_b_0(mesh_5_10_io_in_b_0),
    .io_in_b_1(mesh_5_10_io_in_b_1),
    .io_in_d_0(mesh_5_10_io_in_d_0),
    .io_in_d_1(mesh_5_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_10_io_in_control_1_shift),
    .io_in_id_0(mesh_5_10_io_in_id_0),
    .io_in_id_1(mesh_5_10_io_in_id_1),
    .io_in_last_0(mesh_5_10_io_in_last_0),
    .io_in_last_1(mesh_5_10_io_in_last_1),
    .io_out_a_0(mesh_5_10_io_out_a_0),
    .io_out_a_1(mesh_5_10_io_out_a_1),
    .io_out_c_0(mesh_5_10_io_out_c_0),
    .io_out_c_1(mesh_5_10_io_out_c_1),
    .io_out_b_0(mesh_5_10_io_out_b_0),
    .io_out_b_1(mesh_5_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_10_io_out_control_1_shift),
    .io_out_id_0(mesh_5_10_io_out_id_0),
    .io_out_id_1(mesh_5_10_io_out_id_1),
    .io_out_last_0(mesh_5_10_io_out_last_0),
    .io_out_last_1(mesh_5_10_io_out_last_1),
    .io_in_valid_0(mesh_5_10_io_in_valid_0),
    .io_in_valid_1(mesh_5_10_io_in_valid_1),
    .io_out_valid_0(mesh_5_10_io_out_valid_0),
    .io_out_valid_1(mesh_5_10_io_out_valid_1)
  );
  Tile mesh_5_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_11_clock),
    .io_in_a_0(mesh_5_11_io_in_a_0),
    .io_in_a_1(mesh_5_11_io_in_a_1),
    .io_in_b_0(mesh_5_11_io_in_b_0),
    .io_in_b_1(mesh_5_11_io_in_b_1),
    .io_in_d_0(mesh_5_11_io_in_d_0),
    .io_in_d_1(mesh_5_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_11_io_in_control_1_shift),
    .io_in_id_0(mesh_5_11_io_in_id_0),
    .io_in_id_1(mesh_5_11_io_in_id_1),
    .io_in_last_0(mesh_5_11_io_in_last_0),
    .io_in_last_1(mesh_5_11_io_in_last_1),
    .io_out_a_0(mesh_5_11_io_out_a_0),
    .io_out_a_1(mesh_5_11_io_out_a_1),
    .io_out_c_0(mesh_5_11_io_out_c_0),
    .io_out_c_1(mesh_5_11_io_out_c_1),
    .io_out_b_0(mesh_5_11_io_out_b_0),
    .io_out_b_1(mesh_5_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_11_io_out_control_1_shift),
    .io_out_id_0(mesh_5_11_io_out_id_0),
    .io_out_id_1(mesh_5_11_io_out_id_1),
    .io_out_last_0(mesh_5_11_io_out_last_0),
    .io_out_last_1(mesh_5_11_io_out_last_1),
    .io_in_valid_0(mesh_5_11_io_in_valid_0),
    .io_in_valid_1(mesh_5_11_io_in_valid_1),
    .io_out_valid_0(mesh_5_11_io_out_valid_0),
    .io_out_valid_1(mesh_5_11_io_out_valid_1)
  );
  Tile mesh_5_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_12_clock),
    .io_in_a_0(mesh_5_12_io_in_a_0),
    .io_in_a_1(mesh_5_12_io_in_a_1),
    .io_in_b_0(mesh_5_12_io_in_b_0),
    .io_in_b_1(mesh_5_12_io_in_b_1),
    .io_in_d_0(mesh_5_12_io_in_d_0),
    .io_in_d_1(mesh_5_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_12_io_in_control_1_shift),
    .io_in_id_0(mesh_5_12_io_in_id_0),
    .io_in_id_1(mesh_5_12_io_in_id_1),
    .io_in_last_0(mesh_5_12_io_in_last_0),
    .io_in_last_1(mesh_5_12_io_in_last_1),
    .io_out_a_0(mesh_5_12_io_out_a_0),
    .io_out_a_1(mesh_5_12_io_out_a_1),
    .io_out_c_0(mesh_5_12_io_out_c_0),
    .io_out_c_1(mesh_5_12_io_out_c_1),
    .io_out_b_0(mesh_5_12_io_out_b_0),
    .io_out_b_1(mesh_5_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_12_io_out_control_1_shift),
    .io_out_id_0(mesh_5_12_io_out_id_0),
    .io_out_id_1(mesh_5_12_io_out_id_1),
    .io_out_last_0(mesh_5_12_io_out_last_0),
    .io_out_last_1(mesh_5_12_io_out_last_1),
    .io_in_valid_0(mesh_5_12_io_in_valid_0),
    .io_in_valid_1(mesh_5_12_io_in_valid_1),
    .io_out_valid_0(mesh_5_12_io_out_valid_0),
    .io_out_valid_1(mesh_5_12_io_out_valid_1)
  );
  Tile mesh_5_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_13_clock),
    .io_in_a_0(mesh_5_13_io_in_a_0),
    .io_in_a_1(mesh_5_13_io_in_a_1),
    .io_in_b_0(mesh_5_13_io_in_b_0),
    .io_in_b_1(mesh_5_13_io_in_b_1),
    .io_in_d_0(mesh_5_13_io_in_d_0),
    .io_in_d_1(mesh_5_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_13_io_in_control_1_shift),
    .io_in_id_0(mesh_5_13_io_in_id_0),
    .io_in_id_1(mesh_5_13_io_in_id_1),
    .io_in_last_0(mesh_5_13_io_in_last_0),
    .io_in_last_1(mesh_5_13_io_in_last_1),
    .io_out_a_0(mesh_5_13_io_out_a_0),
    .io_out_a_1(mesh_5_13_io_out_a_1),
    .io_out_c_0(mesh_5_13_io_out_c_0),
    .io_out_c_1(mesh_5_13_io_out_c_1),
    .io_out_b_0(mesh_5_13_io_out_b_0),
    .io_out_b_1(mesh_5_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_13_io_out_control_1_shift),
    .io_out_id_0(mesh_5_13_io_out_id_0),
    .io_out_id_1(mesh_5_13_io_out_id_1),
    .io_out_last_0(mesh_5_13_io_out_last_0),
    .io_out_last_1(mesh_5_13_io_out_last_1),
    .io_in_valid_0(mesh_5_13_io_in_valid_0),
    .io_in_valid_1(mesh_5_13_io_in_valid_1),
    .io_out_valid_0(mesh_5_13_io_out_valid_0),
    .io_out_valid_1(mesh_5_13_io_out_valid_1)
  );
  Tile mesh_5_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_14_clock),
    .io_in_a_0(mesh_5_14_io_in_a_0),
    .io_in_a_1(mesh_5_14_io_in_a_1),
    .io_in_b_0(mesh_5_14_io_in_b_0),
    .io_in_b_1(mesh_5_14_io_in_b_1),
    .io_in_d_0(mesh_5_14_io_in_d_0),
    .io_in_d_1(mesh_5_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_14_io_in_control_1_shift),
    .io_in_id_0(mesh_5_14_io_in_id_0),
    .io_in_id_1(mesh_5_14_io_in_id_1),
    .io_in_last_0(mesh_5_14_io_in_last_0),
    .io_in_last_1(mesh_5_14_io_in_last_1),
    .io_out_a_0(mesh_5_14_io_out_a_0),
    .io_out_a_1(mesh_5_14_io_out_a_1),
    .io_out_c_0(mesh_5_14_io_out_c_0),
    .io_out_c_1(mesh_5_14_io_out_c_1),
    .io_out_b_0(mesh_5_14_io_out_b_0),
    .io_out_b_1(mesh_5_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_14_io_out_control_1_shift),
    .io_out_id_0(mesh_5_14_io_out_id_0),
    .io_out_id_1(mesh_5_14_io_out_id_1),
    .io_out_last_0(mesh_5_14_io_out_last_0),
    .io_out_last_1(mesh_5_14_io_out_last_1),
    .io_in_valid_0(mesh_5_14_io_in_valid_0),
    .io_in_valid_1(mesh_5_14_io_in_valid_1),
    .io_out_valid_0(mesh_5_14_io_out_valid_0),
    .io_out_valid_1(mesh_5_14_io_out_valid_1)
  );
  Tile mesh_5_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_5_15_clock),
    .io_in_a_0(mesh_5_15_io_in_a_0),
    .io_in_a_1(mesh_5_15_io_in_a_1),
    .io_in_b_0(mesh_5_15_io_in_b_0),
    .io_in_b_1(mesh_5_15_io_in_b_1),
    .io_in_d_0(mesh_5_15_io_in_d_0),
    .io_in_d_1(mesh_5_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_5_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_5_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_5_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_5_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_5_15_io_in_control_1_shift),
    .io_in_id_0(mesh_5_15_io_in_id_0),
    .io_in_id_1(mesh_5_15_io_in_id_1),
    .io_in_last_0(mesh_5_15_io_in_last_0),
    .io_in_last_1(mesh_5_15_io_in_last_1),
    .io_out_a_0(mesh_5_15_io_out_a_0),
    .io_out_a_1(mesh_5_15_io_out_a_1),
    .io_out_c_0(mesh_5_15_io_out_c_0),
    .io_out_c_1(mesh_5_15_io_out_c_1),
    .io_out_b_0(mesh_5_15_io_out_b_0),
    .io_out_b_1(mesh_5_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_5_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_5_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_5_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_5_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_5_15_io_out_control_1_shift),
    .io_out_id_0(mesh_5_15_io_out_id_0),
    .io_out_id_1(mesh_5_15_io_out_id_1),
    .io_out_last_0(mesh_5_15_io_out_last_0),
    .io_out_last_1(mesh_5_15_io_out_last_1),
    .io_in_valid_0(mesh_5_15_io_in_valid_0),
    .io_in_valid_1(mesh_5_15_io_in_valid_1),
    .io_out_valid_0(mesh_5_15_io_out_valid_0),
    .io_out_valid_1(mesh_5_15_io_out_valid_1)
  );
  Tile mesh_6_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_0_clock),
    .io_in_a_0(mesh_6_0_io_in_a_0),
    .io_in_a_1(mesh_6_0_io_in_a_1),
    .io_in_b_0(mesh_6_0_io_in_b_0),
    .io_in_b_1(mesh_6_0_io_in_b_1),
    .io_in_d_0(mesh_6_0_io_in_d_0),
    .io_in_d_1(mesh_6_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_0_io_in_control_1_shift),
    .io_in_id_0(mesh_6_0_io_in_id_0),
    .io_in_id_1(mesh_6_0_io_in_id_1),
    .io_in_last_0(mesh_6_0_io_in_last_0),
    .io_in_last_1(mesh_6_0_io_in_last_1),
    .io_out_a_0(mesh_6_0_io_out_a_0),
    .io_out_a_1(mesh_6_0_io_out_a_1),
    .io_out_c_0(mesh_6_0_io_out_c_0),
    .io_out_c_1(mesh_6_0_io_out_c_1),
    .io_out_b_0(mesh_6_0_io_out_b_0),
    .io_out_b_1(mesh_6_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_0_io_out_control_1_shift),
    .io_out_id_0(mesh_6_0_io_out_id_0),
    .io_out_id_1(mesh_6_0_io_out_id_1),
    .io_out_last_0(mesh_6_0_io_out_last_0),
    .io_out_last_1(mesh_6_0_io_out_last_1),
    .io_in_valid_0(mesh_6_0_io_in_valid_0),
    .io_in_valid_1(mesh_6_0_io_in_valid_1),
    .io_out_valid_0(mesh_6_0_io_out_valid_0),
    .io_out_valid_1(mesh_6_0_io_out_valid_1)
  );
  Tile mesh_6_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_1_clock),
    .io_in_a_0(mesh_6_1_io_in_a_0),
    .io_in_a_1(mesh_6_1_io_in_a_1),
    .io_in_b_0(mesh_6_1_io_in_b_0),
    .io_in_b_1(mesh_6_1_io_in_b_1),
    .io_in_d_0(mesh_6_1_io_in_d_0),
    .io_in_d_1(mesh_6_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_1_io_in_control_1_shift),
    .io_in_id_0(mesh_6_1_io_in_id_0),
    .io_in_id_1(mesh_6_1_io_in_id_1),
    .io_in_last_0(mesh_6_1_io_in_last_0),
    .io_in_last_1(mesh_6_1_io_in_last_1),
    .io_out_a_0(mesh_6_1_io_out_a_0),
    .io_out_a_1(mesh_6_1_io_out_a_1),
    .io_out_c_0(mesh_6_1_io_out_c_0),
    .io_out_c_1(mesh_6_1_io_out_c_1),
    .io_out_b_0(mesh_6_1_io_out_b_0),
    .io_out_b_1(mesh_6_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_1_io_out_control_1_shift),
    .io_out_id_0(mesh_6_1_io_out_id_0),
    .io_out_id_1(mesh_6_1_io_out_id_1),
    .io_out_last_0(mesh_6_1_io_out_last_0),
    .io_out_last_1(mesh_6_1_io_out_last_1),
    .io_in_valid_0(mesh_6_1_io_in_valid_0),
    .io_in_valid_1(mesh_6_1_io_in_valid_1),
    .io_out_valid_0(mesh_6_1_io_out_valid_0),
    .io_out_valid_1(mesh_6_1_io_out_valid_1)
  );
  Tile mesh_6_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_2_clock),
    .io_in_a_0(mesh_6_2_io_in_a_0),
    .io_in_a_1(mesh_6_2_io_in_a_1),
    .io_in_b_0(mesh_6_2_io_in_b_0),
    .io_in_b_1(mesh_6_2_io_in_b_1),
    .io_in_d_0(mesh_6_2_io_in_d_0),
    .io_in_d_1(mesh_6_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_2_io_in_control_1_shift),
    .io_in_id_0(mesh_6_2_io_in_id_0),
    .io_in_id_1(mesh_6_2_io_in_id_1),
    .io_in_last_0(mesh_6_2_io_in_last_0),
    .io_in_last_1(mesh_6_2_io_in_last_1),
    .io_out_a_0(mesh_6_2_io_out_a_0),
    .io_out_a_1(mesh_6_2_io_out_a_1),
    .io_out_c_0(mesh_6_2_io_out_c_0),
    .io_out_c_1(mesh_6_2_io_out_c_1),
    .io_out_b_0(mesh_6_2_io_out_b_0),
    .io_out_b_1(mesh_6_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_2_io_out_control_1_shift),
    .io_out_id_0(mesh_6_2_io_out_id_0),
    .io_out_id_1(mesh_6_2_io_out_id_1),
    .io_out_last_0(mesh_6_2_io_out_last_0),
    .io_out_last_1(mesh_6_2_io_out_last_1),
    .io_in_valid_0(mesh_6_2_io_in_valid_0),
    .io_in_valid_1(mesh_6_2_io_in_valid_1),
    .io_out_valid_0(mesh_6_2_io_out_valid_0),
    .io_out_valid_1(mesh_6_2_io_out_valid_1)
  );
  Tile mesh_6_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_3_clock),
    .io_in_a_0(mesh_6_3_io_in_a_0),
    .io_in_a_1(mesh_6_3_io_in_a_1),
    .io_in_b_0(mesh_6_3_io_in_b_0),
    .io_in_b_1(mesh_6_3_io_in_b_1),
    .io_in_d_0(mesh_6_3_io_in_d_0),
    .io_in_d_1(mesh_6_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_3_io_in_control_1_shift),
    .io_in_id_0(mesh_6_3_io_in_id_0),
    .io_in_id_1(mesh_6_3_io_in_id_1),
    .io_in_last_0(mesh_6_3_io_in_last_0),
    .io_in_last_1(mesh_6_3_io_in_last_1),
    .io_out_a_0(mesh_6_3_io_out_a_0),
    .io_out_a_1(mesh_6_3_io_out_a_1),
    .io_out_c_0(mesh_6_3_io_out_c_0),
    .io_out_c_1(mesh_6_3_io_out_c_1),
    .io_out_b_0(mesh_6_3_io_out_b_0),
    .io_out_b_1(mesh_6_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_3_io_out_control_1_shift),
    .io_out_id_0(mesh_6_3_io_out_id_0),
    .io_out_id_1(mesh_6_3_io_out_id_1),
    .io_out_last_0(mesh_6_3_io_out_last_0),
    .io_out_last_1(mesh_6_3_io_out_last_1),
    .io_in_valid_0(mesh_6_3_io_in_valid_0),
    .io_in_valid_1(mesh_6_3_io_in_valid_1),
    .io_out_valid_0(mesh_6_3_io_out_valid_0),
    .io_out_valid_1(mesh_6_3_io_out_valid_1)
  );
  Tile mesh_6_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_4_clock),
    .io_in_a_0(mesh_6_4_io_in_a_0),
    .io_in_a_1(mesh_6_4_io_in_a_1),
    .io_in_b_0(mesh_6_4_io_in_b_0),
    .io_in_b_1(mesh_6_4_io_in_b_1),
    .io_in_d_0(mesh_6_4_io_in_d_0),
    .io_in_d_1(mesh_6_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_4_io_in_control_1_shift),
    .io_in_id_0(mesh_6_4_io_in_id_0),
    .io_in_id_1(mesh_6_4_io_in_id_1),
    .io_in_last_0(mesh_6_4_io_in_last_0),
    .io_in_last_1(mesh_6_4_io_in_last_1),
    .io_out_a_0(mesh_6_4_io_out_a_0),
    .io_out_a_1(mesh_6_4_io_out_a_1),
    .io_out_c_0(mesh_6_4_io_out_c_0),
    .io_out_c_1(mesh_6_4_io_out_c_1),
    .io_out_b_0(mesh_6_4_io_out_b_0),
    .io_out_b_1(mesh_6_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_4_io_out_control_1_shift),
    .io_out_id_0(mesh_6_4_io_out_id_0),
    .io_out_id_1(mesh_6_4_io_out_id_1),
    .io_out_last_0(mesh_6_4_io_out_last_0),
    .io_out_last_1(mesh_6_4_io_out_last_1),
    .io_in_valid_0(mesh_6_4_io_in_valid_0),
    .io_in_valid_1(mesh_6_4_io_in_valid_1),
    .io_out_valid_0(mesh_6_4_io_out_valid_0),
    .io_out_valid_1(mesh_6_4_io_out_valid_1)
  );
  Tile mesh_6_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_5_clock),
    .io_in_a_0(mesh_6_5_io_in_a_0),
    .io_in_a_1(mesh_6_5_io_in_a_1),
    .io_in_b_0(mesh_6_5_io_in_b_0),
    .io_in_b_1(mesh_6_5_io_in_b_1),
    .io_in_d_0(mesh_6_5_io_in_d_0),
    .io_in_d_1(mesh_6_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_5_io_in_control_1_shift),
    .io_in_id_0(mesh_6_5_io_in_id_0),
    .io_in_id_1(mesh_6_5_io_in_id_1),
    .io_in_last_0(mesh_6_5_io_in_last_0),
    .io_in_last_1(mesh_6_5_io_in_last_1),
    .io_out_a_0(mesh_6_5_io_out_a_0),
    .io_out_a_1(mesh_6_5_io_out_a_1),
    .io_out_c_0(mesh_6_5_io_out_c_0),
    .io_out_c_1(mesh_6_5_io_out_c_1),
    .io_out_b_0(mesh_6_5_io_out_b_0),
    .io_out_b_1(mesh_6_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_5_io_out_control_1_shift),
    .io_out_id_0(mesh_6_5_io_out_id_0),
    .io_out_id_1(mesh_6_5_io_out_id_1),
    .io_out_last_0(mesh_6_5_io_out_last_0),
    .io_out_last_1(mesh_6_5_io_out_last_1),
    .io_in_valid_0(mesh_6_5_io_in_valid_0),
    .io_in_valid_1(mesh_6_5_io_in_valid_1),
    .io_out_valid_0(mesh_6_5_io_out_valid_0),
    .io_out_valid_1(mesh_6_5_io_out_valid_1)
  );
  Tile mesh_6_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_6_clock),
    .io_in_a_0(mesh_6_6_io_in_a_0),
    .io_in_a_1(mesh_6_6_io_in_a_1),
    .io_in_b_0(mesh_6_6_io_in_b_0),
    .io_in_b_1(mesh_6_6_io_in_b_1),
    .io_in_d_0(mesh_6_6_io_in_d_0),
    .io_in_d_1(mesh_6_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_6_io_in_control_1_shift),
    .io_in_id_0(mesh_6_6_io_in_id_0),
    .io_in_id_1(mesh_6_6_io_in_id_1),
    .io_in_last_0(mesh_6_6_io_in_last_0),
    .io_in_last_1(mesh_6_6_io_in_last_1),
    .io_out_a_0(mesh_6_6_io_out_a_0),
    .io_out_a_1(mesh_6_6_io_out_a_1),
    .io_out_c_0(mesh_6_6_io_out_c_0),
    .io_out_c_1(mesh_6_6_io_out_c_1),
    .io_out_b_0(mesh_6_6_io_out_b_0),
    .io_out_b_1(mesh_6_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_6_io_out_control_1_shift),
    .io_out_id_0(mesh_6_6_io_out_id_0),
    .io_out_id_1(mesh_6_6_io_out_id_1),
    .io_out_last_0(mesh_6_6_io_out_last_0),
    .io_out_last_1(mesh_6_6_io_out_last_1),
    .io_in_valid_0(mesh_6_6_io_in_valid_0),
    .io_in_valid_1(mesh_6_6_io_in_valid_1),
    .io_out_valid_0(mesh_6_6_io_out_valid_0),
    .io_out_valid_1(mesh_6_6_io_out_valid_1)
  );
  Tile mesh_6_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_7_clock),
    .io_in_a_0(mesh_6_7_io_in_a_0),
    .io_in_a_1(mesh_6_7_io_in_a_1),
    .io_in_b_0(mesh_6_7_io_in_b_0),
    .io_in_b_1(mesh_6_7_io_in_b_1),
    .io_in_d_0(mesh_6_7_io_in_d_0),
    .io_in_d_1(mesh_6_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_7_io_in_control_1_shift),
    .io_in_id_0(mesh_6_7_io_in_id_0),
    .io_in_id_1(mesh_6_7_io_in_id_1),
    .io_in_last_0(mesh_6_7_io_in_last_0),
    .io_in_last_1(mesh_6_7_io_in_last_1),
    .io_out_a_0(mesh_6_7_io_out_a_0),
    .io_out_a_1(mesh_6_7_io_out_a_1),
    .io_out_c_0(mesh_6_7_io_out_c_0),
    .io_out_c_1(mesh_6_7_io_out_c_1),
    .io_out_b_0(mesh_6_7_io_out_b_0),
    .io_out_b_1(mesh_6_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_7_io_out_control_1_shift),
    .io_out_id_0(mesh_6_7_io_out_id_0),
    .io_out_id_1(mesh_6_7_io_out_id_1),
    .io_out_last_0(mesh_6_7_io_out_last_0),
    .io_out_last_1(mesh_6_7_io_out_last_1),
    .io_in_valid_0(mesh_6_7_io_in_valid_0),
    .io_in_valid_1(mesh_6_7_io_in_valid_1),
    .io_out_valid_0(mesh_6_7_io_out_valid_0),
    .io_out_valid_1(mesh_6_7_io_out_valid_1)
  );
  Tile mesh_6_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_8_clock),
    .io_in_a_0(mesh_6_8_io_in_a_0),
    .io_in_a_1(mesh_6_8_io_in_a_1),
    .io_in_b_0(mesh_6_8_io_in_b_0),
    .io_in_b_1(mesh_6_8_io_in_b_1),
    .io_in_d_0(mesh_6_8_io_in_d_0),
    .io_in_d_1(mesh_6_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_8_io_in_control_1_shift),
    .io_in_id_0(mesh_6_8_io_in_id_0),
    .io_in_id_1(mesh_6_8_io_in_id_1),
    .io_in_last_0(mesh_6_8_io_in_last_0),
    .io_in_last_1(mesh_6_8_io_in_last_1),
    .io_out_a_0(mesh_6_8_io_out_a_0),
    .io_out_a_1(mesh_6_8_io_out_a_1),
    .io_out_c_0(mesh_6_8_io_out_c_0),
    .io_out_c_1(mesh_6_8_io_out_c_1),
    .io_out_b_0(mesh_6_8_io_out_b_0),
    .io_out_b_1(mesh_6_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_8_io_out_control_1_shift),
    .io_out_id_0(mesh_6_8_io_out_id_0),
    .io_out_id_1(mesh_6_8_io_out_id_1),
    .io_out_last_0(mesh_6_8_io_out_last_0),
    .io_out_last_1(mesh_6_8_io_out_last_1),
    .io_in_valid_0(mesh_6_8_io_in_valid_0),
    .io_in_valid_1(mesh_6_8_io_in_valid_1),
    .io_out_valid_0(mesh_6_8_io_out_valid_0),
    .io_out_valid_1(mesh_6_8_io_out_valid_1)
  );
  Tile mesh_6_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_9_clock),
    .io_in_a_0(mesh_6_9_io_in_a_0),
    .io_in_a_1(mesh_6_9_io_in_a_1),
    .io_in_b_0(mesh_6_9_io_in_b_0),
    .io_in_b_1(mesh_6_9_io_in_b_1),
    .io_in_d_0(mesh_6_9_io_in_d_0),
    .io_in_d_1(mesh_6_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_9_io_in_control_1_shift),
    .io_in_id_0(mesh_6_9_io_in_id_0),
    .io_in_id_1(mesh_6_9_io_in_id_1),
    .io_in_last_0(mesh_6_9_io_in_last_0),
    .io_in_last_1(mesh_6_9_io_in_last_1),
    .io_out_a_0(mesh_6_9_io_out_a_0),
    .io_out_a_1(mesh_6_9_io_out_a_1),
    .io_out_c_0(mesh_6_9_io_out_c_0),
    .io_out_c_1(mesh_6_9_io_out_c_1),
    .io_out_b_0(mesh_6_9_io_out_b_0),
    .io_out_b_1(mesh_6_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_9_io_out_control_1_shift),
    .io_out_id_0(mesh_6_9_io_out_id_0),
    .io_out_id_1(mesh_6_9_io_out_id_1),
    .io_out_last_0(mesh_6_9_io_out_last_0),
    .io_out_last_1(mesh_6_9_io_out_last_1),
    .io_in_valid_0(mesh_6_9_io_in_valid_0),
    .io_in_valid_1(mesh_6_9_io_in_valid_1),
    .io_out_valid_0(mesh_6_9_io_out_valid_0),
    .io_out_valid_1(mesh_6_9_io_out_valid_1)
  );
  Tile mesh_6_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_10_clock),
    .io_in_a_0(mesh_6_10_io_in_a_0),
    .io_in_a_1(mesh_6_10_io_in_a_1),
    .io_in_b_0(mesh_6_10_io_in_b_0),
    .io_in_b_1(mesh_6_10_io_in_b_1),
    .io_in_d_0(mesh_6_10_io_in_d_0),
    .io_in_d_1(mesh_6_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_10_io_in_control_1_shift),
    .io_in_id_0(mesh_6_10_io_in_id_0),
    .io_in_id_1(mesh_6_10_io_in_id_1),
    .io_in_last_0(mesh_6_10_io_in_last_0),
    .io_in_last_1(mesh_6_10_io_in_last_1),
    .io_out_a_0(mesh_6_10_io_out_a_0),
    .io_out_a_1(mesh_6_10_io_out_a_1),
    .io_out_c_0(mesh_6_10_io_out_c_0),
    .io_out_c_1(mesh_6_10_io_out_c_1),
    .io_out_b_0(mesh_6_10_io_out_b_0),
    .io_out_b_1(mesh_6_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_10_io_out_control_1_shift),
    .io_out_id_0(mesh_6_10_io_out_id_0),
    .io_out_id_1(mesh_6_10_io_out_id_1),
    .io_out_last_0(mesh_6_10_io_out_last_0),
    .io_out_last_1(mesh_6_10_io_out_last_1),
    .io_in_valid_0(mesh_6_10_io_in_valid_0),
    .io_in_valid_1(mesh_6_10_io_in_valid_1),
    .io_out_valid_0(mesh_6_10_io_out_valid_0),
    .io_out_valid_1(mesh_6_10_io_out_valid_1)
  );
  Tile mesh_6_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_11_clock),
    .io_in_a_0(mesh_6_11_io_in_a_0),
    .io_in_a_1(mesh_6_11_io_in_a_1),
    .io_in_b_0(mesh_6_11_io_in_b_0),
    .io_in_b_1(mesh_6_11_io_in_b_1),
    .io_in_d_0(mesh_6_11_io_in_d_0),
    .io_in_d_1(mesh_6_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_11_io_in_control_1_shift),
    .io_in_id_0(mesh_6_11_io_in_id_0),
    .io_in_id_1(mesh_6_11_io_in_id_1),
    .io_in_last_0(mesh_6_11_io_in_last_0),
    .io_in_last_1(mesh_6_11_io_in_last_1),
    .io_out_a_0(mesh_6_11_io_out_a_0),
    .io_out_a_1(mesh_6_11_io_out_a_1),
    .io_out_c_0(mesh_6_11_io_out_c_0),
    .io_out_c_1(mesh_6_11_io_out_c_1),
    .io_out_b_0(mesh_6_11_io_out_b_0),
    .io_out_b_1(mesh_6_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_11_io_out_control_1_shift),
    .io_out_id_0(mesh_6_11_io_out_id_0),
    .io_out_id_1(mesh_6_11_io_out_id_1),
    .io_out_last_0(mesh_6_11_io_out_last_0),
    .io_out_last_1(mesh_6_11_io_out_last_1),
    .io_in_valid_0(mesh_6_11_io_in_valid_0),
    .io_in_valid_1(mesh_6_11_io_in_valid_1),
    .io_out_valid_0(mesh_6_11_io_out_valid_0),
    .io_out_valid_1(mesh_6_11_io_out_valid_1)
  );
  Tile mesh_6_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_12_clock),
    .io_in_a_0(mesh_6_12_io_in_a_0),
    .io_in_a_1(mesh_6_12_io_in_a_1),
    .io_in_b_0(mesh_6_12_io_in_b_0),
    .io_in_b_1(mesh_6_12_io_in_b_1),
    .io_in_d_0(mesh_6_12_io_in_d_0),
    .io_in_d_1(mesh_6_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_12_io_in_control_1_shift),
    .io_in_id_0(mesh_6_12_io_in_id_0),
    .io_in_id_1(mesh_6_12_io_in_id_1),
    .io_in_last_0(mesh_6_12_io_in_last_0),
    .io_in_last_1(mesh_6_12_io_in_last_1),
    .io_out_a_0(mesh_6_12_io_out_a_0),
    .io_out_a_1(mesh_6_12_io_out_a_1),
    .io_out_c_0(mesh_6_12_io_out_c_0),
    .io_out_c_1(mesh_6_12_io_out_c_1),
    .io_out_b_0(mesh_6_12_io_out_b_0),
    .io_out_b_1(mesh_6_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_12_io_out_control_1_shift),
    .io_out_id_0(mesh_6_12_io_out_id_0),
    .io_out_id_1(mesh_6_12_io_out_id_1),
    .io_out_last_0(mesh_6_12_io_out_last_0),
    .io_out_last_1(mesh_6_12_io_out_last_1),
    .io_in_valid_0(mesh_6_12_io_in_valid_0),
    .io_in_valid_1(mesh_6_12_io_in_valid_1),
    .io_out_valid_0(mesh_6_12_io_out_valid_0),
    .io_out_valid_1(mesh_6_12_io_out_valid_1)
  );
  Tile mesh_6_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_13_clock),
    .io_in_a_0(mesh_6_13_io_in_a_0),
    .io_in_a_1(mesh_6_13_io_in_a_1),
    .io_in_b_0(mesh_6_13_io_in_b_0),
    .io_in_b_1(mesh_6_13_io_in_b_1),
    .io_in_d_0(mesh_6_13_io_in_d_0),
    .io_in_d_1(mesh_6_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_13_io_in_control_1_shift),
    .io_in_id_0(mesh_6_13_io_in_id_0),
    .io_in_id_1(mesh_6_13_io_in_id_1),
    .io_in_last_0(mesh_6_13_io_in_last_0),
    .io_in_last_1(mesh_6_13_io_in_last_1),
    .io_out_a_0(mesh_6_13_io_out_a_0),
    .io_out_a_1(mesh_6_13_io_out_a_1),
    .io_out_c_0(mesh_6_13_io_out_c_0),
    .io_out_c_1(mesh_6_13_io_out_c_1),
    .io_out_b_0(mesh_6_13_io_out_b_0),
    .io_out_b_1(mesh_6_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_13_io_out_control_1_shift),
    .io_out_id_0(mesh_6_13_io_out_id_0),
    .io_out_id_1(mesh_6_13_io_out_id_1),
    .io_out_last_0(mesh_6_13_io_out_last_0),
    .io_out_last_1(mesh_6_13_io_out_last_1),
    .io_in_valid_0(mesh_6_13_io_in_valid_0),
    .io_in_valid_1(mesh_6_13_io_in_valid_1),
    .io_out_valid_0(mesh_6_13_io_out_valid_0),
    .io_out_valid_1(mesh_6_13_io_out_valid_1)
  );
  Tile mesh_6_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_14_clock),
    .io_in_a_0(mesh_6_14_io_in_a_0),
    .io_in_a_1(mesh_6_14_io_in_a_1),
    .io_in_b_0(mesh_6_14_io_in_b_0),
    .io_in_b_1(mesh_6_14_io_in_b_1),
    .io_in_d_0(mesh_6_14_io_in_d_0),
    .io_in_d_1(mesh_6_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_14_io_in_control_1_shift),
    .io_in_id_0(mesh_6_14_io_in_id_0),
    .io_in_id_1(mesh_6_14_io_in_id_1),
    .io_in_last_0(mesh_6_14_io_in_last_0),
    .io_in_last_1(mesh_6_14_io_in_last_1),
    .io_out_a_0(mesh_6_14_io_out_a_0),
    .io_out_a_1(mesh_6_14_io_out_a_1),
    .io_out_c_0(mesh_6_14_io_out_c_0),
    .io_out_c_1(mesh_6_14_io_out_c_1),
    .io_out_b_0(mesh_6_14_io_out_b_0),
    .io_out_b_1(mesh_6_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_14_io_out_control_1_shift),
    .io_out_id_0(mesh_6_14_io_out_id_0),
    .io_out_id_1(mesh_6_14_io_out_id_1),
    .io_out_last_0(mesh_6_14_io_out_last_0),
    .io_out_last_1(mesh_6_14_io_out_last_1),
    .io_in_valid_0(mesh_6_14_io_in_valid_0),
    .io_in_valid_1(mesh_6_14_io_in_valid_1),
    .io_out_valid_0(mesh_6_14_io_out_valid_0),
    .io_out_valid_1(mesh_6_14_io_out_valid_1)
  );
  Tile mesh_6_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_6_15_clock),
    .io_in_a_0(mesh_6_15_io_in_a_0),
    .io_in_a_1(mesh_6_15_io_in_a_1),
    .io_in_b_0(mesh_6_15_io_in_b_0),
    .io_in_b_1(mesh_6_15_io_in_b_1),
    .io_in_d_0(mesh_6_15_io_in_d_0),
    .io_in_d_1(mesh_6_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_6_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_6_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_6_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_6_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_6_15_io_in_control_1_shift),
    .io_in_id_0(mesh_6_15_io_in_id_0),
    .io_in_id_1(mesh_6_15_io_in_id_1),
    .io_in_last_0(mesh_6_15_io_in_last_0),
    .io_in_last_1(mesh_6_15_io_in_last_1),
    .io_out_a_0(mesh_6_15_io_out_a_0),
    .io_out_a_1(mesh_6_15_io_out_a_1),
    .io_out_c_0(mesh_6_15_io_out_c_0),
    .io_out_c_1(mesh_6_15_io_out_c_1),
    .io_out_b_0(mesh_6_15_io_out_b_0),
    .io_out_b_1(mesh_6_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_6_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_6_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_6_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_6_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_6_15_io_out_control_1_shift),
    .io_out_id_0(mesh_6_15_io_out_id_0),
    .io_out_id_1(mesh_6_15_io_out_id_1),
    .io_out_last_0(mesh_6_15_io_out_last_0),
    .io_out_last_1(mesh_6_15_io_out_last_1),
    .io_in_valid_0(mesh_6_15_io_in_valid_0),
    .io_in_valid_1(mesh_6_15_io_in_valid_1),
    .io_out_valid_0(mesh_6_15_io_out_valid_0),
    .io_out_valid_1(mesh_6_15_io_out_valid_1)
  );
  Tile mesh_7_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_0_clock),
    .io_in_a_0(mesh_7_0_io_in_a_0),
    .io_in_a_1(mesh_7_0_io_in_a_1),
    .io_in_b_0(mesh_7_0_io_in_b_0),
    .io_in_b_1(mesh_7_0_io_in_b_1),
    .io_in_d_0(mesh_7_0_io_in_d_0),
    .io_in_d_1(mesh_7_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_0_io_in_control_1_shift),
    .io_in_id_0(mesh_7_0_io_in_id_0),
    .io_in_id_1(mesh_7_0_io_in_id_1),
    .io_in_last_0(mesh_7_0_io_in_last_0),
    .io_in_last_1(mesh_7_0_io_in_last_1),
    .io_out_a_0(mesh_7_0_io_out_a_0),
    .io_out_a_1(mesh_7_0_io_out_a_1),
    .io_out_c_0(mesh_7_0_io_out_c_0),
    .io_out_c_1(mesh_7_0_io_out_c_1),
    .io_out_b_0(mesh_7_0_io_out_b_0),
    .io_out_b_1(mesh_7_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_0_io_out_control_1_shift),
    .io_out_id_0(mesh_7_0_io_out_id_0),
    .io_out_id_1(mesh_7_0_io_out_id_1),
    .io_out_last_0(mesh_7_0_io_out_last_0),
    .io_out_last_1(mesh_7_0_io_out_last_1),
    .io_in_valid_0(mesh_7_0_io_in_valid_0),
    .io_in_valid_1(mesh_7_0_io_in_valid_1),
    .io_out_valid_0(mesh_7_0_io_out_valid_0),
    .io_out_valid_1(mesh_7_0_io_out_valid_1)
  );
  Tile mesh_7_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_1_clock),
    .io_in_a_0(mesh_7_1_io_in_a_0),
    .io_in_a_1(mesh_7_1_io_in_a_1),
    .io_in_b_0(mesh_7_1_io_in_b_0),
    .io_in_b_1(mesh_7_1_io_in_b_1),
    .io_in_d_0(mesh_7_1_io_in_d_0),
    .io_in_d_1(mesh_7_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_1_io_in_control_1_shift),
    .io_in_id_0(mesh_7_1_io_in_id_0),
    .io_in_id_1(mesh_7_1_io_in_id_1),
    .io_in_last_0(mesh_7_1_io_in_last_0),
    .io_in_last_1(mesh_7_1_io_in_last_1),
    .io_out_a_0(mesh_7_1_io_out_a_0),
    .io_out_a_1(mesh_7_1_io_out_a_1),
    .io_out_c_0(mesh_7_1_io_out_c_0),
    .io_out_c_1(mesh_7_1_io_out_c_1),
    .io_out_b_0(mesh_7_1_io_out_b_0),
    .io_out_b_1(mesh_7_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_1_io_out_control_1_shift),
    .io_out_id_0(mesh_7_1_io_out_id_0),
    .io_out_id_1(mesh_7_1_io_out_id_1),
    .io_out_last_0(mesh_7_1_io_out_last_0),
    .io_out_last_1(mesh_7_1_io_out_last_1),
    .io_in_valid_0(mesh_7_1_io_in_valid_0),
    .io_in_valid_1(mesh_7_1_io_in_valid_1),
    .io_out_valid_0(mesh_7_1_io_out_valid_0),
    .io_out_valid_1(mesh_7_1_io_out_valid_1)
  );
  Tile mesh_7_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_2_clock),
    .io_in_a_0(mesh_7_2_io_in_a_0),
    .io_in_a_1(mesh_7_2_io_in_a_1),
    .io_in_b_0(mesh_7_2_io_in_b_0),
    .io_in_b_1(mesh_7_2_io_in_b_1),
    .io_in_d_0(mesh_7_2_io_in_d_0),
    .io_in_d_1(mesh_7_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_2_io_in_control_1_shift),
    .io_in_id_0(mesh_7_2_io_in_id_0),
    .io_in_id_1(mesh_7_2_io_in_id_1),
    .io_in_last_0(mesh_7_2_io_in_last_0),
    .io_in_last_1(mesh_7_2_io_in_last_1),
    .io_out_a_0(mesh_7_2_io_out_a_0),
    .io_out_a_1(mesh_7_2_io_out_a_1),
    .io_out_c_0(mesh_7_2_io_out_c_0),
    .io_out_c_1(mesh_7_2_io_out_c_1),
    .io_out_b_0(mesh_7_2_io_out_b_0),
    .io_out_b_1(mesh_7_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_2_io_out_control_1_shift),
    .io_out_id_0(mesh_7_2_io_out_id_0),
    .io_out_id_1(mesh_7_2_io_out_id_1),
    .io_out_last_0(mesh_7_2_io_out_last_0),
    .io_out_last_1(mesh_7_2_io_out_last_1),
    .io_in_valid_0(mesh_7_2_io_in_valid_0),
    .io_in_valid_1(mesh_7_2_io_in_valid_1),
    .io_out_valid_0(mesh_7_2_io_out_valid_0),
    .io_out_valid_1(mesh_7_2_io_out_valid_1)
  );
  Tile mesh_7_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_3_clock),
    .io_in_a_0(mesh_7_3_io_in_a_0),
    .io_in_a_1(mesh_7_3_io_in_a_1),
    .io_in_b_0(mesh_7_3_io_in_b_0),
    .io_in_b_1(mesh_7_3_io_in_b_1),
    .io_in_d_0(mesh_7_3_io_in_d_0),
    .io_in_d_1(mesh_7_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_3_io_in_control_1_shift),
    .io_in_id_0(mesh_7_3_io_in_id_0),
    .io_in_id_1(mesh_7_3_io_in_id_1),
    .io_in_last_0(mesh_7_3_io_in_last_0),
    .io_in_last_1(mesh_7_3_io_in_last_1),
    .io_out_a_0(mesh_7_3_io_out_a_0),
    .io_out_a_1(mesh_7_3_io_out_a_1),
    .io_out_c_0(mesh_7_3_io_out_c_0),
    .io_out_c_1(mesh_7_3_io_out_c_1),
    .io_out_b_0(mesh_7_3_io_out_b_0),
    .io_out_b_1(mesh_7_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_3_io_out_control_1_shift),
    .io_out_id_0(mesh_7_3_io_out_id_0),
    .io_out_id_1(mesh_7_3_io_out_id_1),
    .io_out_last_0(mesh_7_3_io_out_last_0),
    .io_out_last_1(mesh_7_3_io_out_last_1),
    .io_in_valid_0(mesh_7_3_io_in_valid_0),
    .io_in_valid_1(mesh_7_3_io_in_valid_1),
    .io_out_valid_0(mesh_7_3_io_out_valid_0),
    .io_out_valid_1(mesh_7_3_io_out_valid_1)
  );
  Tile mesh_7_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_4_clock),
    .io_in_a_0(mesh_7_4_io_in_a_0),
    .io_in_a_1(mesh_7_4_io_in_a_1),
    .io_in_b_0(mesh_7_4_io_in_b_0),
    .io_in_b_1(mesh_7_4_io_in_b_1),
    .io_in_d_0(mesh_7_4_io_in_d_0),
    .io_in_d_1(mesh_7_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_4_io_in_control_1_shift),
    .io_in_id_0(mesh_7_4_io_in_id_0),
    .io_in_id_1(mesh_7_4_io_in_id_1),
    .io_in_last_0(mesh_7_4_io_in_last_0),
    .io_in_last_1(mesh_7_4_io_in_last_1),
    .io_out_a_0(mesh_7_4_io_out_a_0),
    .io_out_a_1(mesh_7_4_io_out_a_1),
    .io_out_c_0(mesh_7_4_io_out_c_0),
    .io_out_c_1(mesh_7_4_io_out_c_1),
    .io_out_b_0(mesh_7_4_io_out_b_0),
    .io_out_b_1(mesh_7_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_4_io_out_control_1_shift),
    .io_out_id_0(mesh_7_4_io_out_id_0),
    .io_out_id_1(mesh_7_4_io_out_id_1),
    .io_out_last_0(mesh_7_4_io_out_last_0),
    .io_out_last_1(mesh_7_4_io_out_last_1),
    .io_in_valid_0(mesh_7_4_io_in_valid_0),
    .io_in_valid_1(mesh_7_4_io_in_valid_1),
    .io_out_valid_0(mesh_7_4_io_out_valid_0),
    .io_out_valid_1(mesh_7_4_io_out_valid_1)
  );
  Tile mesh_7_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_5_clock),
    .io_in_a_0(mesh_7_5_io_in_a_0),
    .io_in_a_1(mesh_7_5_io_in_a_1),
    .io_in_b_0(mesh_7_5_io_in_b_0),
    .io_in_b_1(mesh_7_5_io_in_b_1),
    .io_in_d_0(mesh_7_5_io_in_d_0),
    .io_in_d_1(mesh_7_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_5_io_in_control_1_shift),
    .io_in_id_0(mesh_7_5_io_in_id_0),
    .io_in_id_1(mesh_7_5_io_in_id_1),
    .io_in_last_0(mesh_7_5_io_in_last_0),
    .io_in_last_1(mesh_7_5_io_in_last_1),
    .io_out_a_0(mesh_7_5_io_out_a_0),
    .io_out_a_1(mesh_7_5_io_out_a_1),
    .io_out_c_0(mesh_7_5_io_out_c_0),
    .io_out_c_1(mesh_7_5_io_out_c_1),
    .io_out_b_0(mesh_7_5_io_out_b_0),
    .io_out_b_1(mesh_7_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_5_io_out_control_1_shift),
    .io_out_id_0(mesh_7_5_io_out_id_0),
    .io_out_id_1(mesh_7_5_io_out_id_1),
    .io_out_last_0(mesh_7_5_io_out_last_0),
    .io_out_last_1(mesh_7_5_io_out_last_1),
    .io_in_valid_0(mesh_7_5_io_in_valid_0),
    .io_in_valid_1(mesh_7_5_io_in_valid_1),
    .io_out_valid_0(mesh_7_5_io_out_valid_0),
    .io_out_valid_1(mesh_7_5_io_out_valid_1)
  );
  Tile mesh_7_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_6_clock),
    .io_in_a_0(mesh_7_6_io_in_a_0),
    .io_in_a_1(mesh_7_6_io_in_a_1),
    .io_in_b_0(mesh_7_6_io_in_b_0),
    .io_in_b_1(mesh_7_6_io_in_b_1),
    .io_in_d_0(mesh_7_6_io_in_d_0),
    .io_in_d_1(mesh_7_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_6_io_in_control_1_shift),
    .io_in_id_0(mesh_7_6_io_in_id_0),
    .io_in_id_1(mesh_7_6_io_in_id_1),
    .io_in_last_0(mesh_7_6_io_in_last_0),
    .io_in_last_1(mesh_7_6_io_in_last_1),
    .io_out_a_0(mesh_7_6_io_out_a_0),
    .io_out_a_1(mesh_7_6_io_out_a_1),
    .io_out_c_0(mesh_7_6_io_out_c_0),
    .io_out_c_1(mesh_7_6_io_out_c_1),
    .io_out_b_0(mesh_7_6_io_out_b_0),
    .io_out_b_1(mesh_7_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_6_io_out_control_1_shift),
    .io_out_id_0(mesh_7_6_io_out_id_0),
    .io_out_id_1(mesh_7_6_io_out_id_1),
    .io_out_last_0(mesh_7_6_io_out_last_0),
    .io_out_last_1(mesh_7_6_io_out_last_1),
    .io_in_valid_0(mesh_7_6_io_in_valid_0),
    .io_in_valid_1(mesh_7_6_io_in_valid_1),
    .io_out_valid_0(mesh_7_6_io_out_valid_0),
    .io_out_valid_1(mesh_7_6_io_out_valid_1)
  );
  Tile mesh_7_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_7_clock),
    .io_in_a_0(mesh_7_7_io_in_a_0),
    .io_in_a_1(mesh_7_7_io_in_a_1),
    .io_in_b_0(mesh_7_7_io_in_b_0),
    .io_in_b_1(mesh_7_7_io_in_b_1),
    .io_in_d_0(mesh_7_7_io_in_d_0),
    .io_in_d_1(mesh_7_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_7_io_in_control_1_shift),
    .io_in_id_0(mesh_7_7_io_in_id_0),
    .io_in_id_1(mesh_7_7_io_in_id_1),
    .io_in_last_0(mesh_7_7_io_in_last_0),
    .io_in_last_1(mesh_7_7_io_in_last_1),
    .io_out_a_0(mesh_7_7_io_out_a_0),
    .io_out_a_1(mesh_7_7_io_out_a_1),
    .io_out_c_0(mesh_7_7_io_out_c_0),
    .io_out_c_1(mesh_7_7_io_out_c_1),
    .io_out_b_0(mesh_7_7_io_out_b_0),
    .io_out_b_1(mesh_7_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_7_io_out_control_1_shift),
    .io_out_id_0(mesh_7_7_io_out_id_0),
    .io_out_id_1(mesh_7_7_io_out_id_1),
    .io_out_last_0(mesh_7_7_io_out_last_0),
    .io_out_last_1(mesh_7_7_io_out_last_1),
    .io_in_valid_0(mesh_7_7_io_in_valid_0),
    .io_in_valid_1(mesh_7_7_io_in_valid_1),
    .io_out_valid_0(mesh_7_7_io_out_valid_0),
    .io_out_valid_1(mesh_7_7_io_out_valid_1)
  );
  Tile mesh_7_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_8_clock),
    .io_in_a_0(mesh_7_8_io_in_a_0),
    .io_in_a_1(mesh_7_8_io_in_a_1),
    .io_in_b_0(mesh_7_8_io_in_b_0),
    .io_in_b_1(mesh_7_8_io_in_b_1),
    .io_in_d_0(mesh_7_8_io_in_d_0),
    .io_in_d_1(mesh_7_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_8_io_in_control_1_shift),
    .io_in_id_0(mesh_7_8_io_in_id_0),
    .io_in_id_1(mesh_7_8_io_in_id_1),
    .io_in_last_0(mesh_7_8_io_in_last_0),
    .io_in_last_1(mesh_7_8_io_in_last_1),
    .io_out_a_0(mesh_7_8_io_out_a_0),
    .io_out_a_1(mesh_7_8_io_out_a_1),
    .io_out_c_0(mesh_7_8_io_out_c_0),
    .io_out_c_1(mesh_7_8_io_out_c_1),
    .io_out_b_0(mesh_7_8_io_out_b_0),
    .io_out_b_1(mesh_7_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_8_io_out_control_1_shift),
    .io_out_id_0(mesh_7_8_io_out_id_0),
    .io_out_id_1(mesh_7_8_io_out_id_1),
    .io_out_last_0(mesh_7_8_io_out_last_0),
    .io_out_last_1(mesh_7_8_io_out_last_1),
    .io_in_valid_0(mesh_7_8_io_in_valid_0),
    .io_in_valid_1(mesh_7_8_io_in_valid_1),
    .io_out_valid_0(mesh_7_8_io_out_valid_0),
    .io_out_valid_1(mesh_7_8_io_out_valid_1)
  );
  Tile mesh_7_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_9_clock),
    .io_in_a_0(mesh_7_9_io_in_a_0),
    .io_in_a_1(mesh_7_9_io_in_a_1),
    .io_in_b_0(mesh_7_9_io_in_b_0),
    .io_in_b_1(mesh_7_9_io_in_b_1),
    .io_in_d_0(mesh_7_9_io_in_d_0),
    .io_in_d_1(mesh_7_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_9_io_in_control_1_shift),
    .io_in_id_0(mesh_7_9_io_in_id_0),
    .io_in_id_1(mesh_7_9_io_in_id_1),
    .io_in_last_0(mesh_7_9_io_in_last_0),
    .io_in_last_1(mesh_7_9_io_in_last_1),
    .io_out_a_0(mesh_7_9_io_out_a_0),
    .io_out_a_1(mesh_7_9_io_out_a_1),
    .io_out_c_0(mesh_7_9_io_out_c_0),
    .io_out_c_1(mesh_7_9_io_out_c_1),
    .io_out_b_0(mesh_7_9_io_out_b_0),
    .io_out_b_1(mesh_7_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_9_io_out_control_1_shift),
    .io_out_id_0(mesh_7_9_io_out_id_0),
    .io_out_id_1(mesh_7_9_io_out_id_1),
    .io_out_last_0(mesh_7_9_io_out_last_0),
    .io_out_last_1(mesh_7_9_io_out_last_1),
    .io_in_valid_0(mesh_7_9_io_in_valid_0),
    .io_in_valid_1(mesh_7_9_io_in_valid_1),
    .io_out_valid_0(mesh_7_9_io_out_valid_0),
    .io_out_valid_1(mesh_7_9_io_out_valid_1)
  );
  Tile mesh_7_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_10_clock),
    .io_in_a_0(mesh_7_10_io_in_a_0),
    .io_in_a_1(mesh_7_10_io_in_a_1),
    .io_in_b_0(mesh_7_10_io_in_b_0),
    .io_in_b_1(mesh_7_10_io_in_b_1),
    .io_in_d_0(mesh_7_10_io_in_d_0),
    .io_in_d_1(mesh_7_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_10_io_in_control_1_shift),
    .io_in_id_0(mesh_7_10_io_in_id_0),
    .io_in_id_1(mesh_7_10_io_in_id_1),
    .io_in_last_0(mesh_7_10_io_in_last_0),
    .io_in_last_1(mesh_7_10_io_in_last_1),
    .io_out_a_0(mesh_7_10_io_out_a_0),
    .io_out_a_1(mesh_7_10_io_out_a_1),
    .io_out_c_0(mesh_7_10_io_out_c_0),
    .io_out_c_1(mesh_7_10_io_out_c_1),
    .io_out_b_0(mesh_7_10_io_out_b_0),
    .io_out_b_1(mesh_7_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_10_io_out_control_1_shift),
    .io_out_id_0(mesh_7_10_io_out_id_0),
    .io_out_id_1(mesh_7_10_io_out_id_1),
    .io_out_last_0(mesh_7_10_io_out_last_0),
    .io_out_last_1(mesh_7_10_io_out_last_1),
    .io_in_valid_0(mesh_7_10_io_in_valid_0),
    .io_in_valid_1(mesh_7_10_io_in_valid_1),
    .io_out_valid_0(mesh_7_10_io_out_valid_0),
    .io_out_valid_1(mesh_7_10_io_out_valid_1)
  );
  Tile mesh_7_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_11_clock),
    .io_in_a_0(mesh_7_11_io_in_a_0),
    .io_in_a_1(mesh_7_11_io_in_a_1),
    .io_in_b_0(mesh_7_11_io_in_b_0),
    .io_in_b_1(mesh_7_11_io_in_b_1),
    .io_in_d_0(mesh_7_11_io_in_d_0),
    .io_in_d_1(mesh_7_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_11_io_in_control_1_shift),
    .io_in_id_0(mesh_7_11_io_in_id_0),
    .io_in_id_1(mesh_7_11_io_in_id_1),
    .io_in_last_0(mesh_7_11_io_in_last_0),
    .io_in_last_1(mesh_7_11_io_in_last_1),
    .io_out_a_0(mesh_7_11_io_out_a_0),
    .io_out_a_1(mesh_7_11_io_out_a_1),
    .io_out_c_0(mesh_7_11_io_out_c_0),
    .io_out_c_1(mesh_7_11_io_out_c_1),
    .io_out_b_0(mesh_7_11_io_out_b_0),
    .io_out_b_1(mesh_7_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_11_io_out_control_1_shift),
    .io_out_id_0(mesh_7_11_io_out_id_0),
    .io_out_id_1(mesh_7_11_io_out_id_1),
    .io_out_last_0(mesh_7_11_io_out_last_0),
    .io_out_last_1(mesh_7_11_io_out_last_1),
    .io_in_valid_0(mesh_7_11_io_in_valid_0),
    .io_in_valid_1(mesh_7_11_io_in_valid_1),
    .io_out_valid_0(mesh_7_11_io_out_valid_0),
    .io_out_valid_1(mesh_7_11_io_out_valid_1)
  );
  Tile mesh_7_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_12_clock),
    .io_in_a_0(mesh_7_12_io_in_a_0),
    .io_in_a_1(mesh_7_12_io_in_a_1),
    .io_in_b_0(mesh_7_12_io_in_b_0),
    .io_in_b_1(mesh_7_12_io_in_b_1),
    .io_in_d_0(mesh_7_12_io_in_d_0),
    .io_in_d_1(mesh_7_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_12_io_in_control_1_shift),
    .io_in_id_0(mesh_7_12_io_in_id_0),
    .io_in_id_1(mesh_7_12_io_in_id_1),
    .io_in_last_0(mesh_7_12_io_in_last_0),
    .io_in_last_1(mesh_7_12_io_in_last_1),
    .io_out_a_0(mesh_7_12_io_out_a_0),
    .io_out_a_1(mesh_7_12_io_out_a_1),
    .io_out_c_0(mesh_7_12_io_out_c_0),
    .io_out_c_1(mesh_7_12_io_out_c_1),
    .io_out_b_0(mesh_7_12_io_out_b_0),
    .io_out_b_1(mesh_7_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_12_io_out_control_1_shift),
    .io_out_id_0(mesh_7_12_io_out_id_0),
    .io_out_id_1(mesh_7_12_io_out_id_1),
    .io_out_last_0(mesh_7_12_io_out_last_0),
    .io_out_last_1(mesh_7_12_io_out_last_1),
    .io_in_valid_0(mesh_7_12_io_in_valid_0),
    .io_in_valid_1(mesh_7_12_io_in_valid_1),
    .io_out_valid_0(mesh_7_12_io_out_valid_0),
    .io_out_valid_1(mesh_7_12_io_out_valid_1)
  );
  Tile mesh_7_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_13_clock),
    .io_in_a_0(mesh_7_13_io_in_a_0),
    .io_in_a_1(mesh_7_13_io_in_a_1),
    .io_in_b_0(mesh_7_13_io_in_b_0),
    .io_in_b_1(mesh_7_13_io_in_b_1),
    .io_in_d_0(mesh_7_13_io_in_d_0),
    .io_in_d_1(mesh_7_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_13_io_in_control_1_shift),
    .io_in_id_0(mesh_7_13_io_in_id_0),
    .io_in_id_1(mesh_7_13_io_in_id_1),
    .io_in_last_0(mesh_7_13_io_in_last_0),
    .io_in_last_1(mesh_7_13_io_in_last_1),
    .io_out_a_0(mesh_7_13_io_out_a_0),
    .io_out_a_1(mesh_7_13_io_out_a_1),
    .io_out_c_0(mesh_7_13_io_out_c_0),
    .io_out_c_1(mesh_7_13_io_out_c_1),
    .io_out_b_0(mesh_7_13_io_out_b_0),
    .io_out_b_1(mesh_7_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_13_io_out_control_1_shift),
    .io_out_id_0(mesh_7_13_io_out_id_0),
    .io_out_id_1(mesh_7_13_io_out_id_1),
    .io_out_last_0(mesh_7_13_io_out_last_0),
    .io_out_last_1(mesh_7_13_io_out_last_1),
    .io_in_valid_0(mesh_7_13_io_in_valid_0),
    .io_in_valid_1(mesh_7_13_io_in_valid_1),
    .io_out_valid_0(mesh_7_13_io_out_valid_0),
    .io_out_valid_1(mesh_7_13_io_out_valid_1)
  );
  Tile mesh_7_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_14_clock),
    .io_in_a_0(mesh_7_14_io_in_a_0),
    .io_in_a_1(mesh_7_14_io_in_a_1),
    .io_in_b_0(mesh_7_14_io_in_b_0),
    .io_in_b_1(mesh_7_14_io_in_b_1),
    .io_in_d_0(mesh_7_14_io_in_d_0),
    .io_in_d_1(mesh_7_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_14_io_in_control_1_shift),
    .io_in_id_0(mesh_7_14_io_in_id_0),
    .io_in_id_1(mesh_7_14_io_in_id_1),
    .io_in_last_0(mesh_7_14_io_in_last_0),
    .io_in_last_1(mesh_7_14_io_in_last_1),
    .io_out_a_0(mesh_7_14_io_out_a_0),
    .io_out_a_1(mesh_7_14_io_out_a_1),
    .io_out_c_0(mesh_7_14_io_out_c_0),
    .io_out_c_1(mesh_7_14_io_out_c_1),
    .io_out_b_0(mesh_7_14_io_out_b_0),
    .io_out_b_1(mesh_7_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_14_io_out_control_1_shift),
    .io_out_id_0(mesh_7_14_io_out_id_0),
    .io_out_id_1(mesh_7_14_io_out_id_1),
    .io_out_last_0(mesh_7_14_io_out_last_0),
    .io_out_last_1(mesh_7_14_io_out_last_1),
    .io_in_valid_0(mesh_7_14_io_in_valid_0),
    .io_in_valid_1(mesh_7_14_io_in_valid_1),
    .io_out_valid_0(mesh_7_14_io_out_valid_0),
    .io_out_valid_1(mesh_7_14_io_out_valid_1)
  );
  Tile mesh_7_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_7_15_clock),
    .io_in_a_0(mesh_7_15_io_in_a_0),
    .io_in_a_1(mesh_7_15_io_in_a_1),
    .io_in_b_0(mesh_7_15_io_in_b_0),
    .io_in_b_1(mesh_7_15_io_in_b_1),
    .io_in_d_0(mesh_7_15_io_in_d_0),
    .io_in_d_1(mesh_7_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_7_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_7_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_7_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_7_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_7_15_io_in_control_1_shift),
    .io_in_id_0(mesh_7_15_io_in_id_0),
    .io_in_id_1(mesh_7_15_io_in_id_1),
    .io_in_last_0(mesh_7_15_io_in_last_0),
    .io_in_last_1(mesh_7_15_io_in_last_1),
    .io_out_a_0(mesh_7_15_io_out_a_0),
    .io_out_a_1(mesh_7_15_io_out_a_1),
    .io_out_c_0(mesh_7_15_io_out_c_0),
    .io_out_c_1(mesh_7_15_io_out_c_1),
    .io_out_b_0(mesh_7_15_io_out_b_0),
    .io_out_b_1(mesh_7_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_7_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_7_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_7_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_7_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_7_15_io_out_control_1_shift),
    .io_out_id_0(mesh_7_15_io_out_id_0),
    .io_out_id_1(mesh_7_15_io_out_id_1),
    .io_out_last_0(mesh_7_15_io_out_last_0),
    .io_out_last_1(mesh_7_15_io_out_last_1),
    .io_in_valid_0(mesh_7_15_io_in_valid_0),
    .io_in_valid_1(mesh_7_15_io_in_valid_1),
    .io_out_valid_0(mesh_7_15_io_out_valid_0),
    .io_out_valid_1(mesh_7_15_io_out_valid_1)
  );
  Tile mesh_8_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_0_clock),
    .io_in_a_0(mesh_8_0_io_in_a_0),
    .io_in_a_1(mesh_8_0_io_in_a_1),
    .io_in_b_0(mesh_8_0_io_in_b_0),
    .io_in_b_1(mesh_8_0_io_in_b_1),
    .io_in_d_0(mesh_8_0_io_in_d_0),
    .io_in_d_1(mesh_8_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_0_io_in_control_1_shift),
    .io_in_id_0(mesh_8_0_io_in_id_0),
    .io_in_id_1(mesh_8_0_io_in_id_1),
    .io_in_last_0(mesh_8_0_io_in_last_0),
    .io_in_last_1(mesh_8_0_io_in_last_1),
    .io_out_a_0(mesh_8_0_io_out_a_0),
    .io_out_a_1(mesh_8_0_io_out_a_1),
    .io_out_c_0(mesh_8_0_io_out_c_0),
    .io_out_c_1(mesh_8_0_io_out_c_1),
    .io_out_b_0(mesh_8_0_io_out_b_0),
    .io_out_b_1(mesh_8_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_0_io_out_control_1_shift),
    .io_out_id_0(mesh_8_0_io_out_id_0),
    .io_out_id_1(mesh_8_0_io_out_id_1),
    .io_out_last_0(mesh_8_0_io_out_last_0),
    .io_out_last_1(mesh_8_0_io_out_last_1),
    .io_in_valid_0(mesh_8_0_io_in_valid_0),
    .io_in_valid_1(mesh_8_0_io_in_valid_1),
    .io_out_valid_0(mesh_8_0_io_out_valid_0),
    .io_out_valid_1(mesh_8_0_io_out_valid_1)
  );
  Tile mesh_8_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_1_clock),
    .io_in_a_0(mesh_8_1_io_in_a_0),
    .io_in_a_1(mesh_8_1_io_in_a_1),
    .io_in_b_0(mesh_8_1_io_in_b_0),
    .io_in_b_1(mesh_8_1_io_in_b_1),
    .io_in_d_0(mesh_8_1_io_in_d_0),
    .io_in_d_1(mesh_8_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_1_io_in_control_1_shift),
    .io_in_id_0(mesh_8_1_io_in_id_0),
    .io_in_id_1(mesh_8_1_io_in_id_1),
    .io_in_last_0(mesh_8_1_io_in_last_0),
    .io_in_last_1(mesh_8_1_io_in_last_1),
    .io_out_a_0(mesh_8_1_io_out_a_0),
    .io_out_a_1(mesh_8_1_io_out_a_1),
    .io_out_c_0(mesh_8_1_io_out_c_0),
    .io_out_c_1(mesh_8_1_io_out_c_1),
    .io_out_b_0(mesh_8_1_io_out_b_0),
    .io_out_b_1(mesh_8_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_1_io_out_control_1_shift),
    .io_out_id_0(mesh_8_1_io_out_id_0),
    .io_out_id_1(mesh_8_1_io_out_id_1),
    .io_out_last_0(mesh_8_1_io_out_last_0),
    .io_out_last_1(mesh_8_1_io_out_last_1),
    .io_in_valid_0(mesh_8_1_io_in_valid_0),
    .io_in_valid_1(mesh_8_1_io_in_valid_1),
    .io_out_valid_0(mesh_8_1_io_out_valid_0),
    .io_out_valid_1(mesh_8_1_io_out_valid_1)
  );
  Tile mesh_8_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_2_clock),
    .io_in_a_0(mesh_8_2_io_in_a_0),
    .io_in_a_1(mesh_8_2_io_in_a_1),
    .io_in_b_0(mesh_8_2_io_in_b_0),
    .io_in_b_1(mesh_8_2_io_in_b_1),
    .io_in_d_0(mesh_8_2_io_in_d_0),
    .io_in_d_1(mesh_8_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_2_io_in_control_1_shift),
    .io_in_id_0(mesh_8_2_io_in_id_0),
    .io_in_id_1(mesh_8_2_io_in_id_1),
    .io_in_last_0(mesh_8_2_io_in_last_0),
    .io_in_last_1(mesh_8_2_io_in_last_1),
    .io_out_a_0(mesh_8_2_io_out_a_0),
    .io_out_a_1(mesh_8_2_io_out_a_1),
    .io_out_c_0(mesh_8_2_io_out_c_0),
    .io_out_c_1(mesh_8_2_io_out_c_1),
    .io_out_b_0(mesh_8_2_io_out_b_0),
    .io_out_b_1(mesh_8_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_2_io_out_control_1_shift),
    .io_out_id_0(mesh_8_2_io_out_id_0),
    .io_out_id_1(mesh_8_2_io_out_id_1),
    .io_out_last_0(mesh_8_2_io_out_last_0),
    .io_out_last_1(mesh_8_2_io_out_last_1),
    .io_in_valid_0(mesh_8_2_io_in_valid_0),
    .io_in_valid_1(mesh_8_2_io_in_valid_1),
    .io_out_valid_0(mesh_8_2_io_out_valid_0),
    .io_out_valid_1(mesh_8_2_io_out_valid_1)
  );
  Tile mesh_8_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_3_clock),
    .io_in_a_0(mesh_8_3_io_in_a_0),
    .io_in_a_1(mesh_8_3_io_in_a_1),
    .io_in_b_0(mesh_8_3_io_in_b_0),
    .io_in_b_1(mesh_8_3_io_in_b_1),
    .io_in_d_0(mesh_8_3_io_in_d_0),
    .io_in_d_1(mesh_8_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_3_io_in_control_1_shift),
    .io_in_id_0(mesh_8_3_io_in_id_0),
    .io_in_id_1(mesh_8_3_io_in_id_1),
    .io_in_last_0(mesh_8_3_io_in_last_0),
    .io_in_last_1(mesh_8_3_io_in_last_1),
    .io_out_a_0(mesh_8_3_io_out_a_0),
    .io_out_a_1(mesh_8_3_io_out_a_1),
    .io_out_c_0(mesh_8_3_io_out_c_0),
    .io_out_c_1(mesh_8_3_io_out_c_1),
    .io_out_b_0(mesh_8_3_io_out_b_0),
    .io_out_b_1(mesh_8_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_3_io_out_control_1_shift),
    .io_out_id_0(mesh_8_3_io_out_id_0),
    .io_out_id_1(mesh_8_3_io_out_id_1),
    .io_out_last_0(mesh_8_3_io_out_last_0),
    .io_out_last_1(mesh_8_3_io_out_last_1),
    .io_in_valid_0(mesh_8_3_io_in_valid_0),
    .io_in_valid_1(mesh_8_3_io_in_valid_1),
    .io_out_valid_0(mesh_8_3_io_out_valid_0),
    .io_out_valid_1(mesh_8_3_io_out_valid_1)
  );
  Tile mesh_8_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_4_clock),
    .io_in_a_0(mesh_8_4_io_in_a_0),
    .io_in_a_1(mesh_8_4_io_in_a_1),
    .io_in_b_0(mesh_8_4_io_in_b_0),
    .io_in_b_1(mesh_8_4_io_in_b_1),
    .io_in_d_0(mesh_8_4_io_in_d_0),
    .io_in_d_1(mesh_8_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_4_io_in_control_1_shift),
    .io_in_id_0(mesh_8_4_io_in_id_0),
    .io_in_id_1(mesh_8_4_io_in_id_1),
    .io_in_last_0(mesh_8_4_io_in_last_0),
    .io_in_last_1(mesh_8_4_io_in_last_1),
    .io_out_a_0(mesh_8_4_io_out_a_0),
    .io_out_a_1(mesh_8_4_io_out_a_1),
    .io_out_c_0(mesh_8_4_io_out_c_0),
    .io_out_c_1(mesh_8_4_io_out_c_1),
    .io_out_b_0(mesh_8_4_io_out_b_0),
    .io_out_b_1(mesh_8_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_4_io_out_control_1_shift),
    .io_out_id_0(mesh_8_4_io_out_id_0),
    .io_out_id_1(mesh_8_4_io_out_id_1),
    .io_out_last_0(mesh_8_4_io_out_last_0),
    .io_out_last_1(mesh_8_4_io_out_last_1),
    .io_in_valid_0(mesh_8_4_io_in_valid_0),
    .io_in_valid_1(mesh_8_4_io_in_valid_1),
    .io_out_valid_0(mesh_8_4_io_out_valid_0),
    .io_out_valid_1(mesh_8_4_io_out_valid_1)
  );
  Tile mesh_8_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_5_clock),
    .io_in_a_0(mesh_8_5_io_in_a_0),
    .io_in_a_1(mesh_8_5_io_in_a_1),
    .io_in_b_0(mesh_8_5_io_in_b_0),
    .io_in_b_1(mesh_8_5_io_in_b_1),
    .io_in_d_0(mesh_8_5_io_in_d_0),
    .io_in_d_1(mesh_8_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_5_io_in_control_1_shift),
    .io_in_id_0(mesh_8_5_io_in_id_0),
    .io_in_id_1(mesh_8_5_io_in_id_1),
    .io_in_last_0(mesh_8_5_io_in_last_0),
    .io_in_last_1(mesh_8_5_io_in_last_1),
    .io_out_a_0(mesh_8_5_io_out_a_0),
    .io_out_a_1(mesh_8_5_io_out_a_1),
    .io_out_c_0(mesh_8_5_io_out_c_0),
    .io_out_c_1(mesh_8_5_io_out_c_1),
    .io_out_b_0(mesh_8_5_io_out_b_0),
    .io_out_b_1(mesh_8_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_5_io_out_control_1_shift),
    .io_out_id_0(mesh_8_5_io_out_id_0),
    .io_out_id_1(mesh_8_5_io_out_id_1),
    .io_out_last_0(mesh_8_5_io_out_last_0),
    .io_out_last_1(mesh_8_5_io_out_last_1),
    .io_in_valid_0(mesh_8_5_io_in_valid_0),
    .io_in_valid_1(mesh_8_5_io_in_valid_1),
    .io_out_valid_0(mesh_8_5_io_out_valid_0),
    .io_out_valid_1(mesh_8_5_io_out_valid_1)
  );
  Tile mesh_8_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_6_clock),
    .io_in_a_0(mesh_8_6_io_in_a_0),
    .io_in_a_1(mesh_8_6_io_in_a_1),
    .io_in_b_0(mesh_8_6_io_in_b_0),
    .io_in_b_1(mesh_8_6_io_in_b_1),
    .io_in_d_0(mesh_8_6_io_in_d_0),
    .io_in_d_1(mesh_8_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_6_io_in_control_1_shift),
    .io_in_id_0(mesh_8_6_io_in_id_0),
    .io_in_id_1(mesh_8_6_io_in_id_1),
    .io_in_last_0(mesh_8_6_io_in_last_0),
    .io_in_last_1(mesh_8_6_io_in_last_1),
    .io_out_a_0(mesh_8_6_io_out_a_0),
    .io_out_a_1(mesh_8_6_io_out_a_1),
    .io_out_c_0(mesh_8_6_io_out_c_0),
    .io_out_c_1(mesh_8_6_io_out_c_1),
    .io_out_b_0(mesh_8_6_io_out_b_0),
    .io_out_b_1(mesh_8_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_6_io_out_control_1_shift),
    .io_out_id_0(mesh_8_6_io_out_id_0),
    .io_out_id_1(mesh_8_6_io_out_id_1),
    .io_out_last_0(mesh_8_6_io_out_last_0),
    .io_out_last_1(mesh_8_6_io_out_last_1),
    .io_in_valid_0(mesh_8_6_io_in_valid_0),
    .io_in_valid_1(mesh_8_6_io_in_valid_1),
    .io_out_valid_0(mesh_8_6_io_out_valid_0),
    .io_out_valid_1(mesh_8_6_io_out_valid_1)
  );
  Tile mesh_8_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_7_clock),
    .io_in_a_0(mesh_8_7_io_in_a_0),
    .io_in_a_1(mesh_8_7_io_in_a_1),
    .io_in_b_0(mesh_8_7_io_in_b_0),
    .io_in_b_1(mesh_8_7_io_in_b_1),
    .io_in_d_0(mesh_8_7_io_in_d_0),
    .io_in_d_1(mesh_8_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_7_io_in_control_1_shift),
    .io_in_id_0(mesh_8_7_io_in_id_0),
    .io_in_id_1(mesh_8_7_io_in_id_1),
    .io_in_last_0(mesh_8_7_io_in_last_0),
    .io_in_last_1(mesh_8_7_io_in_last_1),
    .io_out_a_0(mesh_8_7_io_out_a_0),
    .io_out_a_1(mesh_8_7_io_out_a_1),
    .io_out_c_0(mesh_8_7_io_out_c_0),
    .io_out_c_1(mesh_8_7_io_out_c_1),
    .io_out_b_0(mesh_8_7_io_out_b_0),
    .io_out_b_1(mesh_8_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_7_io_out_control_1_shift),
    .io_out_id_0(mesh_8_7_io_out_id_0),
    .io_out_id_1(mesh_8_7_io_out_id_1),
    .io_out_last_0(mesh_8_7_io_out_last_0),
    .io_out_last_1(mesh_8_7_io_out_last_1),
    .io_in_valid_0(mesh_8_7_io_in_valid_0),
    .io_in_valid_1(mesh_8_7_io_in_valid_1),
    .io_out_valid_0(mesh_8_7_io_out_valid_0),
    .io_out_valid_1(mesh_8_7_io_out_valid_1)
  );
  Tile mesh_8_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_8_clock),
    .io_in_a_0(mesh_8_8_io_in_a_0),
    .io_in_a_1(mesh_8_8_io_in_a_1),
    .io_in_b_0(mesh_8_8_io_in_b_0),
    .io_in_b_1(mesh_8_8_io_in_b_1),
    .io_in_d_0(mesh_8_8_io_in_d_0),
    .io_in_d_1(mesh_8_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_8_io_in_control_1_shift),
    .io_in_id_0(mesh_8_8_io_in_id_0),
    .io_in_id_1(mesh_8_8_io_in_id_1),
    .io_in_last_0(mesh_8_8_io_in_last_0),
    .io_in_last_1(mesh_8_8_io_in_last_1),
    .io_out_a_0(mesh_8_8_io_out_a_0),
    .io_out_a_1(mesh_8_8_io_out_a_1),
    .io_out_c_0(mesh_8_8_io_out_c_0),
    .io_out_c_1(mesh_8_8_io_out_c_1),
    .io_out_b_0(mesh_8_8_io_out_b_0),
    .io_out_b_1(mesh_8_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_8_io_out_control_1_shift),
    .io_out_id_0(mesh_8_8_io_out_id_0),
    .io_out_id_1(mesh_8_8_io_out_id_1),
    .io_out_last_0(mesh_8_8_io_out_last_0),
    .io_out_last_1(mesh_8_8_io_out_last_1),
    .io_in_valid_0(mesh_8_8_io_in_valid_0),
    .io_in_valid_1(mesh_8_8_io_in_valid_1),
    .io_out_valid_0(mesh_8_8_io_out_valid_0),
    .io_out_valid_1(mesh_8_8_io_out_valid_1)
  );
  Tile mesh_8_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_9_clock),
    .io_in_a_0(mesh_8_9_io_in_a_0),
    .io_in_a_1(mesh_8_9_io_in_a_1),
    .io_in_b_0(mesh_8_9_io_in_b_0),
    .io_in_b_1(mesh_8_9_io_in_b_1),
    .io_in_d_0(mesh_8_9_io_in_d_0),
    .io_in_d_1(mesh_8_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_9_io_in_control_1_shift),
    .io_in_id_0(mesh_8_9_io_in_id_0),
    .io_in_id_1(mesh_8_9_io_in_id_1),
    .io_in_last_0(mesh_8_9_io_in_last_0),
    .io_in_last_1(mesh_8_9_io_in_last_1),
    .io_out_a_0(mesh_8_9_io_out_a_0),
    .io_out_a_1(mesh_8_9_io_out_a_1),
    .io_out_c_0(mesh_8_9_io_out_c_0),
    .io_out_c_1(mesh_8_9_io_out_c_1),
    .io_out_b_0(mesh_8_9_io_out_b_0),
    .io_out_b_1(mesh_8_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_9_io_out_control_1_shift),
    .io_out_id_0(mesh_8_9_io_out_id_0),
    .io_out_id_1(mesh_8_9_io_out_id_1),
    .io_out_last_0(mesh_8_9_io_out_last_0),
    .io_out_last_1(mesh_8_9_io_out_last_1),
    .io_in_valid_0(mesh_8_9_io_in_valid_0),
    .io_in_valid_1(mesh_8_9_io_in_valid_1),
    .io_out_valid_0(mesh_8_9_io_out_valid_0),
    .io_out_valid_1(mesh_8_9_io_out_valid_1)
  );
  Tile mesh_8_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_10_clock),
    .io_in_a_0(mesh_8_10_io_in_a_0),
    .io_in_a_1(mesh_8_10_io_in_a_1),
    .io_in_b_0(mesh_8_10_io_in_b_0),
    .io_in_b_1(mesh_8_10_io_in_b_1),
    .io_in_d_0(mesh_8_10_io_in_d_0),
    .io_in_d_1(mesh_8_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_10_io_in_control_1_shift),
    .io_in_id_0(mesh_8_10_io_in_id_0),
    .io_in_id_1(mesh_8_10_io_in_id_1),
    .io_in_last_0(mesh_8_10_io_in_last_0),
    .io_in_last_1(mesh_8_10_io_in_last_1),
    .io_out_a_0(mesh_8_10_io_out_a_0),
    .io_out_a_1(mesh_8_10_io_out_a_1),
    .io_out_c_0(mesh_8_10_io_out_c_0),
    .io_out_c_1(mesh_8_10_io_out_c_1),
    .io_out_b_0(mesh_8_10_io_out_b_0),
    .io_out_b_1(mesh_8_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_10_io_out_control_1_shift),
    .io_out_id_0(mesh_8_10_io_out_id_0),
    .io_out_id_1(mesh_8_10_io_out_id_1),
    .io_out_last_0(mesh_8_10_io_out_last_0),
    .io_out_last_1(mesh_8_10_io_out_last_1),
    .io_in_valid_0(mesh_8_10_io_in_valid_0),
    .io_in_valid_1(mesh_8_10_io_in_valid_1),
    .io_out_valid_0(mesh_8_10_io_out_valid_0),
    .io_out_valid_1(mesh_8_10_io_out_valid_1)
  );
  Tile mesh_8_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_11_clock),
    .io_in_a_0(mesh_8_11_io_in_a_0),
    .io_in_a_1(mesh_8_11_io_in_a_1),
    .io_in_b_0(mesh_8_11_io_in_b_0),
    .io_in_b_1(mesh_8_11_io_in_b_1),
    .io_in_d_0(mesh_8_11_io_in_d_0),
    .io_in_d_1(mesh_8_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_11_io_in_control_1_shift),
    .io_in_id_0(mesh_8_11_io_in_id_0),
    .io_in_id_1(mesh_8_11_io_in_id_1),
    .io_in_last_0(mesh_8_11_io_in_last_0),
    .io_in_last_1(mesh_8_11_io_in_last_1),
    .io_out_a_0(mesh_8_11_io_out_a_0),
    .io_out_a_1(mesh_8_11_io_out_a_1),
    .io_out_c_0(mesh_8_11_io_out_c_0),
    .io_out_c_1(mesh_8_11_io_out_c_1),
    .io_out_b_0(mesh_8_11_io_out_b_0),
    .io_out_b_1(mesh_8_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_11_io_out_control_1_shift),
    .io_out_id_0(mesh_8_11_io_out_id_0),
    .io_out_id_1(mesh_8_11_io_out_id_1),
    .io_out_last_0(mesh_8_11_io_out_last_0),
    .io_out_last_1(mesh_8_11_io_out_last_1),
    .io_in_valid_0(mesh_8_11_io_in_valid_0),
    .io_in_valid_1(mesh_8_11_io_in_valid_1),
    .io_out_valid_0(mesh_8_11_io_out_valid_0),
    .io_out_valid_1(mesh_8_11_io_out_valid_1)
  );
  Tile mesh_8_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_12_clock),
    .io_in_a_0(mesh_8_12_io_in_a_0),
    .io_in_a_1(mesh_8_12_io_in_a_1),
    .io_in_b_0(mesh_8_12_io_in_b_0),
    .io_in_b_1(mesh_8_12_io_in_b_1),
    .io_in_d_0(mesh_8_12_io_in_d_0),
    .io_in_d_1(mesh_8_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_12_io_in_control_1_shift),
    .io_in_id_0(mesh_8_12_io_in_id_0),
    .io_in_id_1(mesh_8_12_io_in_id_1),
    .io_in_last_0(mesh_8_12_io_in_last_0),
    .io_in_last_1(mesh_8_12_io_in_last_1),
    .io_out_a_0(mesh_8_12_io_out_a_0),
    .io_out_a_1(mesh_8_12_io_out_a_1),
    .io_out_c_0(mesh_8_12_io_out_c_0),
    .io_out_c_1(mesh_8_12_io_out_c_1),
    .io_out_b_0(mesh_8_12_io_out_b_0),
    .io_out_b_1(mesh_8_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_12_io_out_control_1_shift),
    .io_out_id_0(mesh_8_12_io_out_id_0),
    .io_out_id_1(mesh_8_12_io_out_id_1),
    .io_out_last_0(mesh_8_12_io_out_last_0),
    .io_out_last_1(mesh_8_12_io_out_last_1),
    .io_in_valid_0(mesh_8_12_io_in_valid_0),
    .io_in_valid_1(mesh_8_12_io_in_valid_1),
    .io_out_valid_0(mesh_8_12_io_out_valid_0),
    .io_out_valid_1(mesh_8_12_io_out_valid_1)
  );
  Tile mesh_8_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_13_clock),
    .io_in_a_0(mesh_8_13_io_in_a_0),
    .io_in_a_1(mesh_8_13_io_in_a_1),
    .io_in_b_0(mesh_8_13_io_in_b_0),
    .io_in_b_1(mesh_8_13_io_in_b_1),
    .io_in_d_0(mesh_8_13_io_in_d_0),
    .io_in_d_1(mesh_8_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_13_io_in_control_1_shift),
    .io_in_id_0(mesh_8_13_io_in_id_0),
    .io_in_id_1(mesh_8_13_io_in_id_1),
    .io_in_last_0(mesh_8_13_io_in_last_0),
    .io_in_last_1(mesh_8_13_io_in_last_1),
    .io_out_a_0(mesh_8_13_io_out_a_0),
    .io_out_a_1(mesh_8_13_io_out_a_1),
    .io_out_c_0(mesh_8_13_io_out_c_0),
    .io_out_c_1(mesh_8_13_io_out_c_1),
    .io_out_b_0(mesh_8_13_io_out_b_0),
    .io_out_b_1(mesh_8_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_13_io_out_control_1_shift),
    .io_out_id_0(mesh_8_13_io_out_id_0),
    .io_out_id_1(mesh_8_13_io_out_id_1),
    .io_out_last_0(mesh_8_13_io_out_last_0),
    .io_out_last_1(mesh_8_13_io_out_last_1),
    .io_in_valid_0(mesh_8_13_io_in_valid_0),
    .io_in_valid_1(mesh_8_13_io_in_valid_1),
    .io_out_valid_0(mesh_8_13_io_out_valid_0),
    .io_out_valid_1(mesh_8_13_io_out_valid_1)
  );
  Tile mesh_8_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_14_clock),
    .io_in_a_0(mesh_8_14_io_in_a_0),
    .io_in_a_1(mesh_8_14_io_in_a_1),
    .io_in_b_0(mesh_8_14_io_in_b_0),
    .io_in_b_1(mesh_8_14_io_in_b_1),
    .io_in_d_0(mesh_8_14_io_in_d_0),
    .io_in_d_1(mesh_8_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_14_io_in_control_1_shift),
    .io_in_id_0(mesh_8_14_io_in_id_0),
    .io_in_id_1(mesh_8_14_io_in_id_1),
    .io_in_last_0(mesh_8_14_io_in_last_0),
    .io_in_last_1(mesh_8_14_io_in_last_1),
    .io_out_a_0(mesh_8_14_io_out_a_0),
    .io_out_a_1(mesh_8_14_io_out_a_1),
    .io_out_c_0(mesh_8_14_io_out_c_0),
    .io_out_c_1(mesh_8_14_io_out_c_1),
    .io_out_b_0(mesh_8_14_io_out_b_0),
    .io_out_b_1(mesh_8_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_14_io_out_control_1_shift),
    .io_out_id_0(mesh_8_14_io_out_id_0),
    .io_out_id_1(mesh_8_14_io_out_id_1),
    .io_out_last_0(mesh_8_14_io_out_last_0),
    .io_out_last_1(mesh_8_14_io_out_last_1),
    .io_in_valid_0(mesh_8_14_io_in_valid_0),
    .io_in_valid_1(mesh_8_14_io_in_valid_1),
    .io_out_valid_0(mesh_8_14_io_out_valid_0),
    .io_out_valid_1(mesh_8_14_io_out_valid_1)
  );
  Tile mesh_8_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_8_15_clock),
    .io_in_a_0(mesh_8_15_io_in_a_0),
    .io_in_a_1(mesh_8_15_io_in_a_1),
    .io_in_b_0(mesh_8_15_io_in_b_0),
    .io_in_b_1(mesh_8_15_io_in_b_1),
    .io_in_d_0(mesh_8_15_io_in_d_0),
    .io_in_d_1(mesh_8_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_8_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_8_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_8_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_8_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_8_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_8_15_io_in_control_1_shift),
    .io_in_id_0(mesh_8_15_io_in_id_0),
    .io_in_id_1(mesh_8_15_io_in_id_1),
    .io_in_last_0(mesh_8_15_io_in_last_0),
    .io_in_last_1(mesh_8_15_io_in_last_1),
    .io_out_a_0(mesh_8_15_io_out_a_0),
    .io_out_a_1(mesh_8_15_io_out_a_1),
    .io_out_c_0(mesh_8_15_io_out_c_0),
    .io_out_c_1(mesh_8_15_io_out_c_1),
    .io_out_b_0(mesh_8_15_io_out_b_0),
    .io_out_b_1(mesh_8_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_8_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_8_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_8_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_8_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_8_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_8_15_io_out_control_1_shift),
    .io_out_id_0(mesh_8_15_io_out_id_0),
    .io_out_id_1(mesh_8_15_io_out_id_1),
    .io_out_last_0(mesh_8_15_io_out_last_0),
    .io_out_last_1(mesh_8_15_io_out_last_1),
    .io_in_valid_0(mesh_8_15_io_in_valid_0),
    .io_in_valid_1(mesh_8_15_io_in_valid_1),
    .io_out_valid_0(mesh_8_15_io_out_valid_0),
    .io_out_valid_1(mesh_8_15_io_out_valid_1)
  );
  Tile mesh_9_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_0_clock),
    .io_in_a_0(mesh_9_0_io_in_a_0),
    .io_in_a_1(mesh_9_0_io_in_a_1),
    .io_in_b_0(mesh_9_0_io_in_b_0),
    .io_in_b_1(mesh_9_0_io_in_b_1),
    .io_in_d_0(mesh_9_0_io_in_d_0),
    .io_in_d_1(mesh_9_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_0_io_in_control_1_shift),
    .io_in_id_0(mesh_9_0_io_in_id_0),
    .io_in_id_1(mesh_9_0_io_in_id_1),
    .io_in_last_0(mesh_9_0_io_in_last_0),
    .io_in_last_1(mesh_9_0_io_in_last_1),
    .io_out_a_0(mesh_9_0_io_out_a_0),
    .io_out_a_1(mesh_9_0_io_out_a_1),
    .io_out_c_0(mesh_9_0_io_out_c_0),
    .io_out_c_1(mesh_9_0_io_out_c_1),
    .io_out_b_0(mesh_9_0_io_out_b_0),
    .io_out_b_1(mesh_9_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_0_io_out_control_1_shift),
    .io_out_id_0(mesh_9_0_io_out_id_0),
    .io_out_id_1(mesh_9_0_io_out_id_1),
    .io_out_last_0(mesh_9_0_io_out_last_0),
    .io_out_last_1(mesh_9_0_io_out_last_1),
    .io_in_valid_0(mesh_9_0_io_in_valid_0),
    .io_in_valid_1(mesh_9_0_io_in_valid_1),
    .io_out_valid_0(mesh_9_0_io_out_valid_0),
    .io_out_valid_1(mesh_9_0_io_out_valid_1)
  );
  Tile mesh_9_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_1_clock),
    .io_in_a_0(mesh_9_1_io_in_a_0),
    .io_in_a_1(mesh_9_1_io_in_a_1),
    .io_in_b_0(mesh_9_1_io_in_b_0),
    .io_in_b_1(mesh_9_1_io_in_b_1),
    .io_in_d_0(mesh_9_1_io_in_d_0),
    .io_in_d_1(mesh_9_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_1_io_in_control_1_shift),
    .io_in_id_0(mesh_9_1_io_in_id_0),
    .io_in_id_1(mesh_9_1_io_in_id_1),
    .io_in_last_0(mesh_9_1_io_in_last_0),
    .io_in_last_1(mesh_9_1_io_in_last_1),
    .io_out_a_0(mesh_9_1_io_out_a_0),
    .io_out_a_1(mesh_9_1_io_out_a_1),
    .io_out_c_0(mesh_9_1_io_out_c_0),
    .io_out_c_1(mesh_9_1_io_out_c_1),
    .io_out_b_0(mesh_9_1_io_out_b_0),
    .io_out_b_1(mesh_9_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_1_io_out_control_1_shift),
    .io_out_id_0(mesh_9_1_io_out_id_0),
    .io_out_id_1(mesh_9_1_io_out_id_1),
    .io_out_last_0(mesh_9_1_io_out_last_0),
    .io_out_last_1(mesh_9_1_io_out_last_1),
    .io_in_valid_0(mesh_9_1_io_in_valid_0),
    .io_in_valid_1(mesh_9_1_io_in_valid_1),
    .io_out_valid_0(mesh_9_1_io_out_valid_0),
    .io_out_valid_1(mesh_9_1_io_out_valid_1)
  );
  Tile mesh_9_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_2_clock),
    .io_in_a_0(mesh_9_2_io_in_a_0),
    .io_in_a_1(mesh_9_2_io_in_a_1),
    .io_in_b_0(mesh_9_2_io_in_b_0),
    .io_in_b_1(mesh_9_2_io_in_b_1),
    .io_in_d_0(mesh_9_2_io_in_d_0),
    .io_in_d_1(mesh_9_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_2_io_in_control_1_shift),
    .io_in_id_0(mesh_9_2_io_in_id_0),
    .io_in_id_1(mesh_9_2_io_in_id_1),
    .io_in_last_0(mesh_9_2_io_in_last_0),
    .io_in_last_1(mesh_9_2_io_in_last_1),
    .io_out_a_0(mesh_9_2_io_out_a_0),
    .io_out_a_1(mesh_9_2_io_out_a_1),
    .io_out_c_0(mesh_9_2_io_out_c_0),
    .io_out_c_1(mesh_9_2_io_out_c_1),
    .io_out_b_0(mesh_9_2_io_out_b_0),
    .io_out_b_1(mesh_9_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_2_io_out_control_1_shift),
    .io_out_id_0(mesh_9_2_io_out_id_0),
    .io_out_id_1(mesh_9_2_io_out_id_1),
    .io_out_last_0(mesh_9_2_io_out_last_0),
    .io_out_last_1(mesh_9_2_io_out_last_1),
    .io_in_valid_0(mesh_9_2_io_in_valid_0),
    .io_in_valid_1(mesh_9_2_io_in_valid_1),
    .io_out_valid_0(mesh_9_2_io_out_valid_0),
    .io_out_valid_1(mesh_9_2_io_out_valid_1)
  );
  Tile mesh_9_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_3_clock),
    .io_in_a_0(mesh_9_3_io_in_a_0),
    .io_in_a_1(mesh_9_3_io_in_a_1),
    .io_in_b_0(mesh_9_3_io_in_b_0),
    .io_in_b_1(mesh_9_3_io_in_b_1),
    .io_in_d_0(mesh_9_3_io_in_d_0),
    .io_in_d_1(mesh_9_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_3_io_in_control_1_shift),
    .io_in_id_0(mesh_9_3_io_in_id_0),
    .io_in_id_1(mesh_9_3_io_in_id_1),
    .io_in_last_0(mesh_9_3_io_in_last_0),
    .io_in_last_1(mesh_9_3_io_in_last_1),
    .io_out_a_0(mesh_9_3_io_out_a_0),
    .io_out_a_1(mesh_9_3_io_out_a_1),
    .io_out_c_0(mesh_9_3_io_out_c_0),
    .io_out_c_1(mesh_9_3_io_out_c_1),
    .io_out_b_0(mesh_9_3_io_out_b_0),
    .io_out_b_1(mesh_9_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_3_io_out_control_1_shift),
    .io_out_id_0(mesh_9_3_io_out_id_0),
    .io_out_id_1(mesh_9_3_io_out_id_1),
    .io_out_last_0(mesh_9_3_io_out_last_0),
    .io_out_last_1(mesh_9_3_io_out_last_1),
    .io_in_valid_0(mesh_9_3_io_in_valid_0),
    .io_in_valid_1(mesh_9_3_io_in_valid_1),
    .io_out_valid_0(mesh_9_3_io_out_valid_0),
    .io_out_valid_1(mesh_9_3_io_out_valid_1)
  );
  Tile mesh_9_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_4_clock),
    .io_in_a_0(mesh_9_4_io_in_a_0),
    .io_in_a_1(mesh_9_4_io_in_a_1),
    .io_in_b_0(mesh_9_4_io_in_b_0),
    .io_in_b_1(mesh_9_4_io_in_b_1),
    .io_in_d_0(mesh_9_4_io_in_d_0),
    .io_in_d_1(mesh_9_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_4_io_in_control_1_shift),
    .io_in_id_0(mesh_9_4_io_in_id_0),
    .io_in_id_1(mesh_9_4_io_in_id_1),
    .io_in_last_0(mesh_9_4_io_in_last_0),
    .io_in_last_1(mesh_9_4_io_in_last_1),
    .io_out_a_0(mesh_9_4_io_out_a_0),
    .io_out_a_1(mesh_9_4_io_out_a_1),
    .io_out_c_0(mesh_9_4_io_out_c_0),
    .io_out_c_1(mesh_9_4_io_out_c_1),
    .io_out_b_0(mesh_9_4_io_out_b_0),
    .io_out_b_1(mesh_9_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_4_io_out_control_1_shift),
    .io_out_id_0(mesh_9_4_io_out_id_0),
    .io_out_id_1(mesh_9_4_io_out_id_1),
    .io_out_last_0(mesh_9_4_io_out_last_0),
    .io_out_last_1(mesh_9_4_io_out_last_1),
    .io_in_valid_0(mesh_9_4_io_in_valid_0),
    .io_in_valid_1(mesh_9_4_io_in_valid_1),
    .io_out_valid_0(mesh_9_4_io_out_valid_0),
    .io_out_valid_1(mesh_9_4_io_out_valid_1)
  );
  Tile mesh_9_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_5_clock),
    .io_in_a_0(mesh_9_5_io_in_a_0),
    .io_in_a_1(mesh_9_5_io_in_a_1),
    .io_in_b_0(mesh_9_5_io_in_b_0),
    .io_in_b_1(mesh_9_5_io_in_b_1),
    .io_in_d_0(mesh_9_5_io_in_d_0),
    .io_in_d_1(mesh_9_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_5_io_in_control_1_shift),
    .io_in_id_0(mesh_9_5_io_in_id_0),
    .io_in_id_1(mesh_9_5_io_in_id_1),
    .io_in_last_0(mesh_9_5_io_in_last_0),
    .io_in_last_1(mesh_9_5_io_in_last_1),
    .io_out_a_0(mesh_9_5_io_out_a_0),
    .io_out_a_1(mesh_9_5_io_out_a_1),
    .io_out_c_0(mesh_9_5_io_out_c_0),
    .io_out_c_1(mesh_9_5_io_out_c_1),
    .io_out_b_0(mesh_9_5_io_out_b_0),
    .io_out_b_1(mesh_9_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_5_io_out_control_1_shift),
    .io_out_id_0(mesh_9_5_io_out_id_0),
    .io_out_id_1(mesh_9_5_io_out_id_1),
    .io_out_last_0(mesh_9_5_io_out_last_0),
    .io_out_last_1(mesh_9_5_io_out_last_1),
    .io_in_valid_0(mesh_9_5_io_in_valid_0),
    .io_in_valid_1(mesh_9_5_io_in_valid_1),
    .io_out_valid_0(mesh_9_5_io_out_valid_0),
    .io_out_valid_1(mesh_9_5_io_out_valid_1)
  );
  Tile mesh_9_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_6_clock),
    .io_in_a_0(mesh_9_6_io_in_a_0),
    .io_in_a_1(mesh_9_6_io_in_a_1),
    .io_in_b_0(mesh_9_6_io_in_b_0),
    .io_in_b_1(mesh_9_6_io_in_b_1),
    .io_in_d_0(mesh_9_6_io_in_d_0),
    .io_in_d_1(mesh_9_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_6_io_in_control_1_shift),
    .io_in_id_0(mesh_9_6_io_in_id_0),
    .io_in_id_1(mesh_9_6_io_in_id_1),
    .io_in_last_0(mesh_9_6_io_in_last_0),
    .io_in_last_1(mesh_9_6_io_in_last_1),
    .io_out_a_0(mesh_9_6_io_out_a_0),
    .io_out_a_1(mesh_9_6_io_out_a_1),
    .io_out_c_0(mesh_9_6_io_out_c_0),
    .io_out_c_1(mesh_9_6_io_out_c_1),
    .io_out_b_0(mesh_9_6_io_out_b_0),
    .io_out_b_1(mesh_9_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_6_io_out_control_1_shift),
    .io_out_id_0(mesh_9_6_io_out_id_0),
    .io_out_id_1(mesh_9_6_io_out_id_1),
    .io_out_last_0(mesh_9_6_io_out_last_0),
    .io_out_last_1(mesh_9_6_io_out_last_1),
    .io_in_valid_0(mesh_9_6_io_in_valid_0),
    .io_in_valid_1(mesh_9_6_io_in_valid_1),
    .io_out_valid_0(mesh_9_6_io_out_valid_0),
    .io_out_valid_1(mesh_9_6_io_out_valid_1)
  );
  Tile mesh_9_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_7_clock),
    .io_in_a_0(mesh_9_7_io_in_a_0),
    .io_in_a_1(mesh_9_7_io_in_a_1),
    .io_in_b_0(mesh_9_7_io_in_b_0),
    .io_in_b_1(mesh_9_7_io_in_b_1),
    .io_in_d_0(mesh_9_7_io_in_d_0),
    .io_in_d_1(mesh_9_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_7_io_in_control_1_shift),
    .io_in_id_0(mesh_9_7_io_in_id_0),
    .io_in_id_1(mesh_9_7_io_in_id_1),
    .io_in_last_0(mesh_9_7_io_in_last_0),
    .io_in_last_1(mesh_9_7_io_in_last_1),
    .io_out_a_0(mesh_9_7_io_out_a_0),
    .io_out_a_1(mesh_9_7_io_out_a_1),
    .io_out_c_0(mesh_9_7_io_out_c_0),
    .io_out_c_1(mesh_9_7_io_out_c_1),
    .io_out_b_0(mesh_9_7_io_out_b_0),
    .io_out_b_1(mesh_9_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_7_io_out_control_1_shift),
    .io_out_id_0(mesh_9_7_io_out_id_0),
    .io_out_id_1(mesh_9_7_io_out_id_1),
    .io_out_last_0(mesh_9_7_io_out_last_0),
    .io_out_last_1(mesh_9_7_io_out_last_1),
    .io_in_valid_0(mesh_9_7_io_in_valid_0),
    .io_in_valid_1(mesh_9_7_io_in_valid_1),
    .io_out_valid_0(mesh_9_7_io_out_valid_0),
    .io_out_valid_1(mesh_9_7_io_out_valid_1)
  );
  Tile mesh_9_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_8_clock),
    .io_in_a_0(mesh_9_8_io_in_a_0),
    .io_in_a_1(mesh_9_8_io_in_a_1),
    .io_in_b_0(mesh_9_8_io_in_b_0),
    .io_in_b_1(mesh_9_8_io_in_b_1),
    .io_in_d_0(mesh_9_8_io_in_d_0),
    .io_in_d_1(mesh_9_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_8_io_in_control_1_shift),
    .io_in_id_0(mesh_9_8_io_in_id_0),
    .io_in_id_1(mesh_9_8_io_in_id_1),
    .io_in_last_0(mesh_9_8_io_in_last_0),
    .io_in_last_1(mesh_9_8_io_in_last_1),
    .io_out_a_0(mesh_9_8_io_out_a_0),
    .io_out_a_1(mesh_9_8_io_out_a_1),
    .io_out_c_0(mesh_9_8_io_out_c_0),
    .io_out_c_1(mesh_9_8_io_out_c_1),
    .io_out_b_0(mesh_9_8_io_out_b_0),
    .io_out_b_1(mesh_9_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_8_io_out_control_1_shift),
    .io_out_id_0(mesh_9_8_io_out_id_0),
    .io_out_id_1(mesh_9_8_io_out_id_1),
    .io_out_last_0(mesh_9_8_io_out_last_0),
    .io_out_last_1(mesh_9_8_io_out_last_1),
    .io_in_valid_0(mesh_9_8_io_in_valid_0),
    .io_in_valid_1(mesh_9_8_io_in_valid_1),
    .io_out_valid_0(mesh_9_8_io_out_valid_0),
    .io_out_valid_1(mesh_9_8_io_out_valid_1)
  );
  Tile mesh_9_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_9_clock),
    .io_in_a_0(mesh_9_9_io_in_a_0),
    .io_in_a_1(mesh_9_9_io_in_a_1),
    .io_in_b_0(mesh_9_9_io_in_b_0),
    .io_in_b_1(mesh_9_9_io_in_b_1),
    .io_in_d_0(mesh_9_9_io_in_d_0),
    .io_in_d_1(mesh_9_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_9_io_in_control_1_shift),
    .io_in_id_0(mesh_9_9_io_in_id_0),
    .io_in_id_1(mesh_9_9_io_in_id_1),
    .io_in_last_0(mesh_9_9_io_in_last_0),
    .io_in_last_1(mesh_9_9_io_in_last_1),
    .io_out_a_0(mesh_9_9_io_out_a_0),
    .io_out_a_1(mesh_9_9_io_out_a_1),
    .io_out_c_0(mesh_9_9_io_out_c_0),
    .io_out_c_1(mesh_9_9_io_out_c_1),
    .io_out_b_0(mesh_9_9_io_out_b_0),
    .io_out_b_1(mesh_9_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_9_io_out_control_1_shift),
    .io_out_id_0(mesh_9_9_io_out_id_0),
    .io_out_id_1(mesh_9_9_io_out_id_1),
    .io_out_last_0(mesh_9_9_io_out_last_0),
    .io_out_last_1(mesh_9_9_io_out_last_1),
    .io_in_valid_0(mesh_9_9_io_in_valid_0),
    .io_in_valid_1(mesh_9_9_io_in_valid_1),
    .io_out_valid_0(mesh_9_9_io_out_valid_0),
    .io_out_valid_1(mesh_9_9_io_out_valid_1)
  );
  Tile mesh_9_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_10_clock),
    .io_in_a_0(mesh_9_10_io_in_a_0),
    .io_in_a_1(mesh_9_10_io_in_a_1),
    .io_in_b_0(mesh_9_10_io_in_b_0),
    .io_in_b_1(mesh_9_10_io_in_b_1),
    .io_in_d_0(mesh_9_10_io_in_d_0),
    .io_in_d_1(mesh_9_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_10_io_in_control_1_shift),
    .io_in_id_0(mesh_9_10_io_in_id_0),
    .io_in_id_1(mesh_9_10_io_in_id_1),
    .io_in_last_0(mesh_9_10_io_in_last_0),
    .io_in_last_1(mesh_9_10_io_in_last_1),
    .io_out_a_0(mesh_9_10_io_out_a_0),
    .io_out_a_1(mesh_9_10_io_out_a_1),
    .io_out_c_0(mesh_9_10_io_out_c_0),
    .io_out_c_1(mesh_9_10_io_out_c_1),
    .io_out_b_0(mesh_9_10_io_out_b_0),
    .io_out_b_1(mesh_9_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_10_io_out_control_1_shift),
    .io_out_id_0(mesh_9_10_io_out_id_0),
    .io_out_id_1(mesh_9_10_io_out_id_1),
    .io_out_last_0(mesh_9_10_io_out_last_0),
    .io_out_last_1(mesh_9_10_io_out_last_1),
    .io_in_valid_0(mesh_9_10_io_in_valid_0),
    .io_in_valid_1(mesh_9_10_io_in_valid_1),
    .io_out_valid_0(mesh_9_10_io_out_valid_0),
    .io_out_valid_1(mesh_9_10_io_out_valid_1)
  );
  Tile mesh_9_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_11_clock),
    .io_in_a_0(mesh_9_11_io_in_a_0),
    .io_in_a_1(mesh_9_11_io_in_a_1),
    .io_in_b_0(mesh_9_11_io_in_b_0),
    .io_in_b_1(mesh_9_11_io_in_b_1),
    .io_in_d_0(mesh_9_11_io_in_d_0),
    .io_in_d_1(mesh_9_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_11_io_in_control_1_shift),
    .io_in_id_0(mesh_9_11_io_in_id_0),
    .io_in_id_1(mesh_9_11_io_in_id_1),
    .io_in_last_0(mesh_9_11_io_in_last_0),
    .io_in_last_1(mesh_9_11_io_in_last_1),
    .io_out_a_0(mesh_9_11_io_out_a_0),
    .io_out_a_1(mesh_9_11_io_out_a_1),
    .io_out_c_0(mesh_9_11_io_out_c_0),
    .io_out_c_1(mesh_9_11_io_out_c_1),
    .io_out_b_0(mesh_9_11_io_out_b_0),
    .io_out_b_1(mesh_9_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_11_io_out_control_1_shift),
    .io_out_id_0(mesh_9_11_io_out_id_0),
    .io_out_id_1(mesh_9_11_io_out_id_1),
    .io_out_last_0(mesh_9_11_io_out_last_0),
    .io_out_last_1(mesh_9_11_io_out_last_1),
    .io_in_valid_0(mesh_9_11_io_in_valid_0),
    .io_in_valid_1(mesh_9_11_io_in_valid_1),
    .io_out_valid_0(mesh_9_11_io_out_valid_0),
    .io_out_valid_1(mesh_9_11_io_out_valid_1)
  );
  Tile mesh_9_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_12_clock),
    .io_in_a_0(mesh_9_12_io_in_a_0),
    .io_in_a_1(mesh_9_12_io_in_a_1),
    .io_in_b_0(mesh_9_12_io_in_b_0),
    .io_in_b_1(mesh_9_12_io_in_b_1),
    .io_in_d_0(mesh_9_12_io_in_d_0),
    .io_in_d_1(mesh_9_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_12_io_in_control_1_shift),
    .io_in_id_0(mesh_9_12_io_in_id_0),
    .io_in_id_1(mesh_9_12_io_in_id_1),
    .io_in_last_0(mesh_9_12_io_in_last_0),
    .io_in_last_1(mesh_9_12_io_in_last_1),
    .io_out_a_0(mesh_9_12_io_out_a_0),
    .io_out_a_1(mesh_9_12_io_out_a_1),
    .io_out_c_0(mesh_9_12_io_out_c_0),
    .io_out_c_1(mesh_9_12_io_out_c_1),
    .io_out_b_0(mesh_9_12_io_out_b_0),
    .io_out_b_1(mesh_9_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_12_io_out_control_1_shift),
    .io_out_id_0(mesh_9_12_io_out_id_0),
    .io_out_id_1(mesh_9_12_io_out_id_1),
    .io_out_last_0(mesh_9_12_io_out_last_0),
    .io_out_last_1(mesh_9_12_io_out_last_1),
    .io_in_valid_0(mesh_9_12_io_in_valid_0),
    .io_in_valid_1(mesh_9_12_io_in_valid_1),
    .io_out_valid_0(mesh_9_12_io_out_valid_0),
    .io_out_valid_1(mesh_9_12_io_out_valid_1)
  );
  Tile mesh_9_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_13_clock),
    .io_in_a_0(mesh_9_13_io_in_a_0),
    .io_in_a_1(mesh_9_13_io_in_a_1),
    .io_in_b_0(mesh_9_13_io_in_b_0),
    .io_in_b_1(mesh_9_13_io_in_b_1),
    .io_in_d_0(mesh_9_13_io_in_d_0),
    .io_in_d_1(mesh_9_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_13_io_in_control_1_shift),
    .io_in_id_0(mesh_9_13_io_in_id_0),
    .io_in_id_1(mesh_9_13_io_in_id_1),
    .io_in_last_0(mesh_9_13_io_in_last_0),
    .io_in_last_1(mesh_9_13_io_in_last_1),
    .io_out_a_0(mesh_9_13_io_out_a_0),
    .io_out_a_1(mesh_9_13_io_out_a_1),
    .io_out_c_0(mesh_9_13_io_out_c_0),
    .io_out_c_1(mesh_9_13_io_out_c_1),
    .io_out_b_0(mesh_9_13_io_out_b_0),
    .io_out_b_1(mesh_9_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_13_io_out_control_1_shift),
    .io_out_id_0(mesh_9_13_io_out_id_0),
    .io_out_id_1(mesh_9_13_io_out_id_1),
    .io_out_last_0(mesh_9_13_io_out_last_0),
    .io_out_last_1(mesh_9_13_io_out_last_1),
    .io_in_valid_0(mesh_9_13_io_in_valid_0),
    .io_in_valid_1(mesh_9_13_io_in_valid_1),
    .io_out_valid_0(mesh_9_13_io_out_valid_0),
    .io_out_valid_1(mesh_9_13_io_out_valid_1)
  );
  Tile mesh_9_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_14_clock),
    .io_in_a_0(mesh_9_14_io_in_a_0),
    .io_in_a_1(mesh_9_14_io_in_a_1),
    .io_in_b_0(mesh_9_14_io_in_b_0),
    .io_in_b_1(mesh_9_14_io_in_b_1),
    .io_in_d_0(mesh_9_14_io_in_d_0),
    .io_in_d_1(mesh_9_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_14_io_in_control_1_shift),
    .io_in_id_0(mesh_9_14_io_in_id_0),
    .io_in_id_1(mesh_9_14_io_in_id_1),
    .io_in_last_0(mesh_9_14_io_in_last_0),
    .io_in_last_1(mesh_9_14_io_in_last_1),
    .io_out_a_0(mesh_9_14_io_out_a_0),
    .io_out_a_1(mesh_9_14_io_out_a_1),
    .io_out_c_0(mesh_9_14_io_out_c_0),
    .io_out_c_1(mesh_9_14_io_out_c_1),
    .io_out_b_0(mesh_9_14_io_out_b_0),
    .io_out_b_1(mesh_9_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_14_io_out_control_1_shift),
    .io_out_id_0(mesh_9_14_io_out_id_0),
    .io_out_id_1(mesh_9_14_io_out_id_1),
    .io_out_last_0(mesh_9_14_io_out_last_0),
    .io_out_last_1(mesh_9_14_io_out_last_1),
    .io_in_valid_0(mesh_9_14_io_in_valid_0),
    .io_in_valid_1(mesh_9_14_io_in_valid_1),
    .io_out_valid_0(mesh_9_14_io_out_valid_0),
    .io_out_valid_1(mesh_9_14_io_out_valid_1)
  );
  Tile mesh_9_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_9_15_clock),
    .io_in_a_0(mesh_9_15_io_in_a_0),
    .io_in_a_1(mesh_9_15_io_in_a_1),
    .io_in_b_0(mesh_9_15_io_in_b_0),
    .io_in_b_1(mesh_9_15_io_in_b_1),
    .io_in_d_0(mesh_9_15_io_in_d_0),
    .io_in_d_1(mesh_9_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_9_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_9_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_9_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_9_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_9_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_9_15_io_in_control_1_shift),
    .io_in_id_0(mesh_9_15_io_in_id_0),
    .io_in_id_1(mesh_9_15_io_in_id_1),
    .io_in_last_0(mesh_9_15_io_in_last_0),
    .io_in_last_1(mesh_9_15_io_in_last_1),
    .io_out_a_0(mesh_9_15_io_out_a_0),
    .io_out_a_1(mesh_9_15_io_out_a_1),
    .io_out_c_0(mesh_9_15_io_out_c_0),
    .io_out_c_1(mesh_9_15_io_out_c_1),
    .io_out_b_0(mesh_9_15_io_out_b_0),
    .io_out_b_1(mesh_9_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_9_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_9_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_9_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_9_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_9_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_9_15_io_out_control_1_shift),
    .io_out_id_0(mesh_9_15_io_out_id_0),
    .io_out_id_1(mesh_9_15_io_out_id_1),
    .io_out_last_0(mesh_9_15_io_out_last_0),
    .io_out_last_1(mesh_9_15_io_out_last_1),
    .io_in_valid_0(mesh_9_15_io_in_valid_0),
    .io_in_valid_1(mesh_9_15_io_in_valid_1),
    .io_out_valid_0(mesh_9_15_io_out_valid_0),
    .io_out_valid_1(mesh_9_15_io_out_valid_1)
  );
  Tile mesh_10_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_0_clock),
    .io_in_a_0(mesh_10_0_io_in_a_0),
    .io_in_a_1(mesh_10_0_io_in_a_1),
    .io_in_b_0(mesh_10_0_io_in_b_0),
    .io_in_b_1(mesh_10_0_io_in_b_1),
    .io_in_d_0(mesh_10_0_io_in_d_0),
    .io_in_d_1(mesh_10_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_0_io_in_control_1_shift),
    .io_in_id_0(mesh_10_0_io_in_id_0),
    .io_in_id_1(mesh_10_0_io_in_id_1),
    .io_in_last_0(mesh_10_0_io_in_last_0),
    .io_in_last_1(mesh_10_0_io_in_last_1),
    .io_out_a_0(mesh_10_0_io_out_a_0),
    .io_out_a_1(mesh_10_0_io_out_a_1),
    .io_out_c_0(mesh_10_0_io_out_c_0),
    .io_out_c_1(mesh_10_0_io_out_c_1),
    .io_out_b_0(mesh_10_0_io_out_b_0),
    .io_out_b_1(mesh_10_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_0_io_out_control_1_shift),
    .io_out_id_0(mesh_10_0_io_out_id_0),
    .io_out_id_1(mesh_10_0_io_out_id_1),
    .io_out_last_0(mesh_10_0_io_out_last_0),
    .io_out_last_1(mesh_10_0_io_out_last_1),
    .io_in_valid_0(mesh_10_0_io_in_valid_0),
    .io_in_valid_1(mesh_10_0_io_in_valid_1),
    .io_out_valid_0(mesh_10_0_io_out_valid_0),
    .io_out_valid_1(mesh_10_0_io_out_valid_1)
  );
  Tile mesh_10_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_1_clock),
    .io_in_a_0(mesh_10_1_io_in_a_0),
    .io_in_a_1(mesh_10_1_io_in_a_1),
    .io_in_b_0(mesh_10_1_io_in_b_0),
    .io_in_b_1(mesh_10_1_io_in_b_1),
    .io_in_d_0(mesh_10_1_io_in_d_0),
    .io_in_d_1(mesh_10_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_1_io_in_control_1_shift),
    .io_in_id_0(mesh_10_1_io_in_id_0),
    .io_in_id_1(mesh_10_1_io_in_id_1),
    .io_in_last_0(mesh_10_1_io_in_last_0),
    .io_in_last_1(mesh_10_1_io_in_last_1),
    .io_out_a_0(mesh_10_1_io_out_a_0),
    .io_out_a_1(mesh_10_1_io_out_a_1),
    .io_out_c_0(mesh_10_1_io_out_c_0),
    .io_out_c_1(mesh_10_1_io_out_c_1),
    .io_out_b_0(mesh_10_1_io_out_b_0),
    .io_out_b_1(mesh_10_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_1_io_out_control_1_shift),
    .io_out_id_0(mesh_10_1_io_out_id_0),
    .io_out_id_1(mesh_10_1_io_out_id_1),
    .io_out_last_0(mesh_10_1_io_out_last_0),
    .io_out_last_1(mesh_10_1_io_out_last_1),
    .io_in_valid_0(mesh_10_1_io_in_valid_0),
    .io_in_valid_1(mesh_10_1_io_in_valid_1),
    .io_out_valid_0(mesh_10_1_io_out_valid_0),
    .io_out_valid_1(mesh_10_1_io_out_valid_1)
  );
  Tile mesh_10_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_2_clock),
    .io_in_a_0(mesh_10_2_io_in_a_0),
    .io_in_a_1(mesh_10_2_io_in_a_1),
    .io_in_b_0(mesh_10_2_io_in_b_0),
    .io_in_b_1(mesh_10_2_io_in_b_1),
    .io_in_d_0(mesh_10_2_io_in_d_0),
    .io_in_d_1(mesh_10_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_2_io_in_control_1_shift),
    .io_in_id_0(mesh_10_2_io_in_id_0),
    .io_in_id_1(mesh_10_2_io_in_id_1),
    .io_in_last_0(mesh_10_2_io_in_last_0),
    .io_in_last_1(mesh_10_2_io_in_last_1),
    .io_out_a_0(mesh_10_2_io_out_a_0),
    .io_out_a_1(mesh_10_2_io_out_a_1),
    .io_out_c_0(mesh_10_2_io_out_c_0),
    .io_out_c_1(mesh_10_2_io_out_c_1),
    .io_out_b_0(mesh_10_2_io_out_b_0),
    .io_out_b_1(mesh_10_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_2_io_out_control_1_shift),
    .io_out_id_0(mesh_10_2_io_out_id_0),
    .io_out_id_1(mesh_10_2_io_out_id_1),
    .io_out_last_0(mesh_10_2_io_out_last_0),
    .io_out_last_1(mesh_10_2_io_out_last_1),
    .io_in_valid_0(mesh_10_2_io_in_valid_0),
    .io_in_valid_1(mesh_10_2_io_in_valid_1),
    .io_out_valid_0(mesh_10_2_io_out_valid_0),
    .io_out_valid_1(mesh_10_2_io_out_valid_1)
  );
  Tile mesh_10_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_3_clock),
    .io_in_a_0(mesh_10_3_io_in_a_0),
    .io_in_a_1(mesh_10_3_io_in_a_1),
    .io_in_b_0(mesh_10_3_io_in_b_0),
    .io_in_b_1(mesh_10_3_io_in_b_1),
    .io_in_d_0(mesh_10_3_io_in_d_0),
    .io_in_d_1(mesh_10_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_3_io_in_control_1_shift),
    .io_in_id_0(mesh_10_3_io_in_id_0),
    .io_in_id_1(mesh_10_3_io_in_id_1),
    .io_in_last_0(mesh_10_3_io_in_last_0),
    .io_in_last_1(mesh_10_3_io_in_last_1),
    .io_out_a_0(mesh_10_3_io_out_a_0),
    .io_out_a_1(mesh_10_3_io_out_a_1),
    .io_out_c_0(mesh_10_3_io_out_c_0),
    .io_out_c_1(mesh_10_3_io_out_c_1),
    .io_out_b_0(mesh_10_3_io_out_b_0),
    .io_out_b_1(mesh_10_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_3_io_out_control_1_shift),
    .io_out_id_0(mesh_10_3_io_out_id_0),
    .io_out_id_1(mesh_10_3_io_out_id_1),
    .io_out_last_0(mesh_10_3_io_out_last_0),
    .io_out_last_1(mesh_10_3_io_out_last_1),
    .io_in_valid_0(mesh_10_3_io_in_valid_0),
    .io_in_valid_1(mesh_10_3_io_in_valid_1),
    .io_out_valid_0(mesh_10_3_io_out_valid_0),
    .io_out_valid_1(mesh_10_3_io_out_valid_1)
  );
  Tile mesh_10_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_4_clock),
    .io_in_a_0(mesh_10_4_io_in_a_0),
    .io_in_a_1(mesh_10_4_io_in_a_1),
    .io_in_b_0(mesh_10_4_io_in_b_0),
    .io_in_b_1(mesh_10_4_io_in_b_1),
    .io_in_d_0(mesh_10_4_io_in_d_0),
    .io_in_d_1(mesh_10_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_4_io_in_control_1_shift),
    .io_in_id_0(mesh_10_4_io_in_id_0),
    .io_in_id_1(mesh_10_4_io_in_id_1),
    .io_in_last_0(mesh_10_4_io_in_last_0),
    .io_in_last_1(mesh_10_4_io_in_last_1),
    .io_out_a_0(mesh_10_4_io_out_a_0),
    .io_out_a_1(mesh_10_4_io_out_a_1),
    .io_out_c_0(mesh_10_4_io_out_c_0),
    .io_out_c_1(mesh_10_4_io_out_c_1),
    .io_out_b_0(mesh_10_4_io_out_b_0),
    .io_out_b_1(mesh_10_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_4_io_out_control_1_shift),
    .io_out_id_0(mesh_10_4_io_out_id_0),
    .io_out_id_1(mesh_10_4_io_out_id_1),
    .io_out_last_0(mesh_10_4_io_out_last_0),
    .io_out_last_1(mesh_10_4_io_out_last_1),
    .io_in_valid_0(mesh_10_4_io_in_valid_0),
    .io_in_valid_1(mesh_10_4_io_in_valid_1),
    .io_out_valid_0(mesh_10_4_io_out_valid_0),
    .io_out_valid_1(mesh_10_4_io_out_valid_1)
  );
  Tile mesh_10_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_5_clock),
    .io_in_a_0(mesh_10_5_io_in_a_0),
    .io_in_a_1(mesh_10_5_io_in_a_1),
    .io_in_b_0(mesh_10_5_io_in_b_0),
    .io_in_b_1(mesh_10_5_io_in_b_1),
    .io_in_d_0(mesh_10_5_io_in_d_0),
    .io_in_d_1(mesh_10_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_5_io_in_control_1_shift),
    .io_in_id_0(mesh_10_5_io_in_id_0),
    .io_in_id_1(mesh_10_5_io_in_id_1),
    .io_in_last_0(mesh_10_5_io_in_last_0),
    .io_in_last_1(mesh_10_5_io_in_last_1),
    .io_out_a_0(mesh_10_5_io_out_a_0),
    .io_out_a_1(mesh_10_5_io_out_a_1),
    .io_out_c_0(mesh_10_5_io_out_c_0),
    .io_out_c_1(mesh_10_5_io_out_c_1),
    .io_out_b_0(mesh_10_5_io_out_b_0),
    .io_out_b_1(mesh_10_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_5_io_out_control_1_shift),
    .io_out_id_0(mesh_10_5_io_out_id_0),
    .io_out_id_1(mesh_10_5_io_out_id_1),
    .io_out_last_0(mesh_10_5_io_out_last_0),
    .io_out_last_1(mesh_10_5_io_out_last_1),
    .io_in_valid_0(mesh_10_5_io_in_valid_0),
    .io_in_valid_1(mesh_10_5_io_in_valid_1),
    .io_out_valid_0(mesh_10_5_io_out_valid_0),
    .io_out_valid_1(mesh_10_5_io_out_valid_1)
  );
  Tile mesh_10_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_6_clock),
    .io_in_a_0(mesh_10_6_io_in_a_0),
    .io_in_a_1(mesh_10_6_io_in_a_1),
    .io_in_b_0(mesh_10_6_io_in_b_0),
    .io_in_b_1(mesh_10_6_io_in_b_1),
    .io_in_d_0(mesh_10_6_io_in_d_0),
    .io_in_d_1(mesh_10_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_6_io_in_control_1_shift),
    .io_in_id_0(mesh_10_6_io_in_id_0),
    .io_in_id_1(mesh_10_6_io_in_id_1),
    .io_in_last_0(mesh_10_6_io_in_last_0),
    .io_in_last_1(mesh_10_6_io_in_last_1),
    .io_out_a_0(mesh_10_6_io_out_a_0),
    .io_out_a_1(mesh_10_6_io_out_a_1),
    .io_out_c_0(mesh_10_6_io_out_c_0),
    .io_out_c_1(mesh_10_6_io_out_c_1),
    .io_out_b_0(mesh_10_6_io_out_b_0),
    .io_out_b_1(mesh_10_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_6_io_out_control_1_shift),
    .io_out_id_0(mesh_10_6_io_out_id_0),
    .io_out_id_1(mesh_10_6_io_out_id_1),
    .io_out_last_0(mesh_10_6_io_out_last_0),
    .io_out_last_1(mesh_10_6_io_out_last_1),
    .io_in_valid_0(mesh_10_6_io_in_valid_0),
    .io_in_valid_1(mesh_10_6_io_in_valid_1),
    .io_out_valid_0(mesh_10_6_io_out_valid_0),
    .io_out_valid_1(mesh_10_6_io_out_valid_1)
  );
  Tile mesh_10_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_7_clock),
    .io_in_a_0(mesh_10_7_io_in_a_0),
    .io_in_a_1(mesh_10_7_io_in_a_1),
    .io_in_b_0(mesh_10_7_io_in_b_0),
    .io_in_b_1(mesh_10_7_io_in_b_1),
    .io_in_d_0(mesh_10_7_io_in_d_0),
    .io_in_d_1(mesh_10_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_7_io_in_control_1_shift),
    .io_in_id_0(mesh_10_7_io_in_id_0),
    .io_in_id_1(mesh_10_7_io_in_id_1),
    .io_in_last_0(mesh_10_7_io_in_last_0),
    .io_in_last_1(mesh_10_7_io_in_last_1),
    .io_out_a_0(mesh_10_7_io_out_a_0),
    .io_out_a_1(mesh_10_7_io_out_a_1),
    .io_out_c_0(mesh_10_7_io_out_c_0),
    .io_out_c_1(mesh_10_7_io_out_c_1),
    .io_out_b_0(mesh_10_7_io_out_b_0),
    .io_out_b_1(mesh_10_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_7_io_out_control_1_shift),
    .io_out_id_0(mesh_10_7_io_out_id_0),
    .io_out_id_1(mesh_10_7_io_out_id_1),
    .io_out_last_0(mesh_10_7_io_out_last_0),
    .io_out_last_1(mesh_10_7_io_out_last_1),
    .io_in_valid_0(mesh_10_7_io_in_valid_0),
    .io_in_valid_1(mesh_10_7_io_in_valid_1),
    .io_out_valid_0(mesh_10_7_io_out_valid_0),
    .io_out_valid_1(mesh_10_7_io_out_valid_1)
  );
  Tile mesh_10_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_8_clock),
    .io_in_a_0(mesh_10_8_io_in_a_0),
    .io_in_a_1(mesh_10_8_io_in_a_1),
    .io_in_b_0(mesh_10_8_io_in_b_0),
    .io_in_b_1(mesh_10_8_io_in_b_1),
    .io_in_d_0(mesh_10_8_io_in_d_0),
    .io_in_d_1(mesh_10_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_8_io_in_control_1_shift),
    .io_in_id_0(mesh_10_8_io_in_id_0),
    .io_in_id_1(mesh_10_8_io_in_id_1),
    .io_in_last_0(mesh_10_8_io_in_last_0),
    .io_in_last_1(mesh_10_8_io_in_last_1),
    .io_out_a_0(mesh_10_8_io_out_a_0),
    .io_out_a_1(mesh_10_8_io_out_a_1),
    .io_out_c_0(mesh_10_8_io_out_c_0),
    .io_out_c_1(mesh_10_8_io_out_c_1),
    .io_out_b_0(mesh_10_8_io_out_b_0),
    .io_out_b_1(mesh_10_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_8_io_out_control_1_shift),
    .io_out_id_0(mesh_10_8_io_out_id_0),
    .io_out_id_1(mesh_10_8_io_out_id_1),
    .io_out_last_0(mesh_10_8_io_out_last_0),
    .io_out_last_1(mesh_10_8_io_out_last_1),
    .io_in_valid_0(mesh_10_8_io_in_valid_0),
    .io_in_valid_1(mesh_10_8_io_in_valid_1),
    .io_out_valid_0(mesh_10_8_io_out_valid_0),
    .io_out_valid_1(mesh_10_8_io_out_valid_1)
  );
  Tile mesh_10_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_9_clock),
    .io_in_a_0(mesh_10_9_io_in_a_0),
    .io_in_a_1(mesh_10_9_io_in_a_1),
    .io_in_b_0(mesh_10_9_io_in_b_0),
    .io_in_b_1(mesh_10_9_io_in_b_1),
    .io_in_d_0(mesh_10_9_io_in_d_0),
    .io_in_d_1(mesh_10_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_9_io_in_control_1_shift),
    .io_in_id_0(mesh_10_9_io_in_id_0),
    .io_in_id_1(mesh_10_9_io_in_id_1),
    .io_in_last_0(mesh_10_9_io_in_last_0),
    .io_in_last_1(mesh_10_9_io_in_last_1),
    .io_out_a_0(mesh_10_9_io_out_a_0),
    .io_out_a_1(mesh_10_9_io_out_a_1),
    .io_out_c_0(mesh_10_9_io_out_c_0),
    .io_out_c_1(mesh_10_9_io_out_c_1),
    .io_out_b_0(mesh_10_9_io_out_b_0),
    .io_out_b_1(mesh_10_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_9_io_out_control_1_shift),
    .io_out_id_0(mesh_10_9_io_out_id_0),
    .io_out_id_1(mesh_10_9_io_out_id_1),
    .io_out_last_0(mesh_10_9_io_out_last_0),
    .io_out_last_1(mesh_10_9_io_out_last_1),
    .io_in_valid_0(mesh_10_9_io_in_valid_0),
    .io_in_valid_1(mesh_10_9_io_in_valid_1),
    .io_out_valid_0(mesh_10_9_io_out_valid_0),
    .io_out_valid_1(mesh_10_9_io_out_valid_1)
  );
  Tile mesh_10_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_10_clock),
    .io_in_a_0(mesh_10_10_io_in_a_0),
    .io_in_a_1(mesh_10_10_io_in_a_1),
    .io_in_b_0(mesh_10_10_io_in_b_0),
    .io_in_b_1(mesh_10_10_io_in_b_1),
    .io_in_d_0(mesh_10_10_io_in_d_0),
    .io_in_d_1(mesh_10_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_10_io_in_control_1_shift),
    .io_in_id_0(mesh_10_10_io_in_id_0),
    .io_in_id_1(mesh_10_10_io_in_id_1),
    .io_in_last_0(mesh_10_10_io_in_last_0),
    .io_in_last_1(mesh_10_10_io_in_last_1),
    .io_out_a_0(mesh_10_10_io_out_a_0),
    .io_out_a_1(mesh_10_10_io_out_a_1),
    .io_out_c_0(mesh_10_10_io_out_c_0),
    .io_out_c_1(mesh_10_10_io_out_c_1),
    .io_out_b_0(mesh_10_10_io_out_b_0),
    .io_out_b_1(mesh_10_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_10_io_out_control_1_shift),
    .io_out_id_0(mesh_10_10_io_out_id_0),
    .io_out_id_1(mesh_10_10_io_out_id_1),
    .io_out_last_0(mesh_10_10_io_out_last_0),
    .io_out_last_1(mesh_10_10_io_out_last_1),
    .io_in_valid_0(mesh_10_10_io_in_valid_0),
    .io_in_valid_1(mesh_10_10_io_in_valid_1),
    .io_out_valid_0(mesh_10_10_io_out_valid_0),
    .io_out_valid_1(mesh_10_10_io_out_valid_1)
  );
  Tile mesh_10_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_11_clock),
    .io_in_a_0(mesh_10_11_io_in_a_0),
    .io_in_a_1(mesh_10_11_io_in_a_1),
    .io_in_b_0(mesh_10_11_io_in_b_0),
    .io_in_b_1(mesh_10_11_io_in_b_1),
    .io_in_d_0(mesh_10_11_io_in_d_0),
    .io_in_d_1(mesh_10_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_11_io_in_control_1_shift),
    .io_in_id_0(mesh_10_11_io_in_id_0),
    .io_in_id_1(mesh_10_11_io_in_id_1),
    .io_in_last_0(mesh_10_11_io_in_last_0),
    .io_in_last_1(mesh_10_11_io_in_last_1),
    .io_out_a_0(mesh_10_11_io_out_a_0),
    .io_out_a_1(mesh_10_11_io_out_a_1),
    .io_out_c_0(mesh_10_11_io_out_c_0),
    .io_out_c_1(mesh_10_11_io_out_c_1),
    .io_out_b_0(mesh_10_11_io_out_b_0),
    .io_out_b_1(mesh_10_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_11_io_out_control_1_shift),
    .io_out_id_0(mesh_10_11_io_out_id_0),
    .io_out_id_1(mesh_10_11_io_out_id_1),
    .io_out_last_0(mesh_10_11_io_out_last_0),
    .io_out_last_1(mesh_10_11_io_out_last_1),
    .io_in_valid_0(mesh_10_11_io_in_valid_0),
    .io_in_valid_1(mesh_10_11_io_in_valid_1),
    .io_out_valid_0(mesh_10_11_io_out_valid_0),
    .io_out_valid_1(mesh_10_11_io_out_valid_1)
  );
  Tile mesh_10_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_12_clock),
    .io_in_a_0(mesh_10_12_io_in_a_0),
    .io_in_a_1(mesh_10_12_io_in_a_1),
    .io_in_b_0(mesh_10_12_io_in_b_0),
    .io_in_b_1(mesh_10_12_io_in_b_1),
    .io_in_d_0(mesh_10_12_io_in_d_0),
    .io_in_d_1(mesh_10_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_12_io_in_control_1_shift),
    .io_in_id_0(mesh_10_12_io_in_id_0),
    .io_in_id_1(mesh_10_12_io_in_id_1),
    .io_in_last_0(mesh_10_12_io_in_last_0),
    .io_in_last_1(mesh_10_12_io_in_last_1),
    .io_out_a_0(mesh_10_12_io_out_a_0),
    .io_out_a_1(mesh_10_12_io_out_a_1),
    .io_out_c_0(mesh_10_12_io_out_c_0),
    .io_out_c_1(mesh_10_12_io_out_c_1),
    .io_out_b_0(mesh_10_12_io_out_b_0),
    .io_out_b_1(mesh_10_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_12_io_out_control_1_shift),
    .io_out_id_0(mesh_10_12_io_out_id_0),
    .io_out_id_1(mesh_10_12_io_out_id_1),
    .io_out_last_0(mesh_10_12_io_out_last_0),
    .io_out_last_1(mesh_10_12_io_out_last_1),
    .io_in_valid_0(mesh_10_12_io_in_valid_0),
    .io_in_valid_1(mesh_10_12_io_in_valid_1),
    .io_out_valid_0(mesh_10_12_io_out_valid_0),
    .io_out_valid_1(mesh_10_12_io_out_valid_1)
  );
  Tile mesh_10_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_13_clock),
    .io_in_a_0(mesh_10_13_io_in_a_0),
    .io_in_a_1(mesh_10_13_io_in_a_1),
    .io_in_b_0(mesh_10_13_io_in_b_0),
    .io_in_b_1(mesh_10_13_io_in_b_1),
    .io_in_d_0(mesh_10_13_io_in_d_0),
    .io_in_d_1(mesh_10_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_13_io_in_control_1_shift),
    .io_in_id_0(mesh_10_13_io_in_id_0),
    .io_in_id_1(mesh_10_13_io_in_id_1),
    .io_in_last_0(mesh_10_13_io_in_last_0),
    .io_in_last_1(mesh_10_13_io_in_last_1),
    .io_out_a_0(mesh_10_13_io_out_a_0),
    .io_out_a_1(mesh_10_13_io_out_a_1),
    .io_out_c_0(mesh_10_13_io_out_c_0),
    .io_out_c_1(mesh_10_13_io_out_c_1),
    .io_out_b_0(mesh_10_13_io_out_b_0),
    .io_out_b_1(mesh_10_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_13_io_out_control_1_shift),
    .io_out_id_0(mesh_10_13_io_out_id_0),
    .io_out_id_1(mesh_10_13_io_out_id_1),
    .io_out_last_0(mesh_10_13_io_out_last_0),
    .io_out_last_1(mesh_10_13_io_out_last_1),
    .io_in_valid_0(mesh_10_13_io_in_valid_0),
    .io_in_valid_1(mesh_10_13_io_in_valid_1),
    .io_out_valid_0(mesh_10_13_io_out_valid_0),
    .io_out_valid_1(mesh_10_13_io_out_valid_1)
  );
  Tile mesh_10_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_14_clock),
    .io_in_a_0(mesh_10_14_io_in_a_0),
    .io_in_a_1(mesh_10_14_io_in_a_1),
    .io_in_b_0(mesh_10_14_io_in_b_0),
    .io_in_b_1(mesh_10_14_io_in_b_1),
    .io_in_d_0(mesh_10_14_io_in_d_0),
    .io_in_d_1(mesh_10_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_14_io_in_control_1_shift),
    .io_in_id_0(mesh_10_14_io_in_id_0),
    .io_in_id_1(mesh_10_14_io_in_id_1),
    .io_in_last_0(mesh_10_14_io_in_last_0),
    .io_in_last_1(mesh_10_14_io_in_last_1),
    .io_out_a_0(mesh_10_14_io_out_a_0),
    .io_out_a_1(mesh_10_14_io_out_a_1),
    .io_out_c_0(mesh_10_14_io_out_c_0),
    .io_out_c_1(mesh_10_14_io_out_c_1),
    .io_out_b_0(mesh_10_14_io_out_b_0),
    .io_out_b_1(mesh_10_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_14_io_out_control_1_shift),
    .io_out_id_0(mesh_10_14_io_out_id_0),
    .io_out_id_1(mesh_10_14_io_out_id_1),
    .io_out_last_0(mesh_10_14_io_out_last_0),
    .io_out_last_1(mesh_10_14_io_out_last_1),
    .io_in_valid_0(mesh_10_14_io_in_valid_0),
    .io_in_valid_1(mesh_10_14_io_in_valid_1),
    .io_out_valid_0(mesh_10_14_io_out_valid_0),
    .io_out_valid_1(mesh_10_14_io_out_valid_1)
  );
  Tile mesh_10_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_10_15_clock),
    .io_in_a_0(mesh_10_15_io_in_a_0),
    .io_in_a_1(mesh_10_15_io_in_a_1),
    .io_in_b_0(mesh_10_15_io_in_b_0),
    .io_in_b_1(mesh_10_15_io_in_b_1),
    .io_in_d_0(mesh_10_15_io_in_d_0),
    .io_in_d_1(mesh_10_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_10_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_10_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_10_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_10_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_10_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_10_15_io_in_control_1_shift),
    .io_in_id_0(mesh_10_15_io_in_id_0),
    .io_in_id_1(mesh_10_15_io_in_id_1),
    .io_in_last_0(mesh_10_15_io_in_last_0),
    .io_in_last_1(mesh_10_15_io_in_last_1),
    .io_out_a_0(mesh_10_15_io_out_a_0),
    .io_out_a_1(mesh_10_15_io_out_a_1),
    .io_out_c_0(mesh_10_15_io_out_c_0),
    .io_out_c_1(mesh_10_15_io_out_c_1),
    .io_out_b_0(mesh_10_15_io_out_b_0),
    .io_out_b_1(mesh_10_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_10_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_10_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_10_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_10_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_10_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_10_15_io_out_control_1_shift),
    .io_out_id_0(mesh_10_15_io_out_id_0),
    .io_out_id_1(mesh_10_15_io_out_id_1),
    .io_out_last_0(mesh_10_15_io_out_last_0),
    .io_out_last_1(mesh_10_15_io_out_last_1),
    .io_in_valid_0(mesh_10_15_io_in_valid_0),
    .io_in_valid_1(mesh_10_15_io_in_valid_1),
    .io_out_valid_0(mesh_10_15_io_out_valid_0),
    .io_out_valid_1(mesh_10_15_io_out_valid_1)
  );
  Tile mesh_11_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_0_clock),
    .io_in_a_0(mesh_11_0_io_in_a_0),
    .io_in_a_1(mesh_11_0_io_in_a_1),
    .io_in_b_0(mesh_11_0_io_in_b_0),
    .io_in_b_1(mesh_11_0_io_in_b_1),
    .io_in_d_0(mesh_11_0_io_in_d_0),
    .io_in_d_1(mesh_11_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_0_io_in_control_1_shift),
    .io_in_id_0(mesh_11_0_io_in_id_0),
    .io_in_id_1(mesh_11_0_io_in_id_1),
    .io_in_last_0(mesh_11_0_io_in_last_0),
    .io_in_last_1(mesh_11_0_io_in_last_1),
    .io_out_a_0(mesh_11_0_io_out_a_0),
    .io_out_a_1(mesh_11_0_io_out_a_1),
    .io_out_c_0(mesh_11_0_io_out_c_0),
    .io_out_c_1(mesh_11_0_io_out_c_1),
    .io_out_b_0(mesh_11_0_io_out_b_0),
    .io_out_b_1(mesh_11_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_0_io_out_control_1_shift),
    .io_out_id_0(mesh_11_0_io_out_id_0),
    .io_out_id_1(mesh_11_0_io_out_id_1),
    .io_out_last_0(mesh_11_0_io_out_last_0),
    .io_out_last_1(mesh_11_0_io_out_last_1),
    .io_in_valid_0(mesh_11_0_io_in_valid_0),
    .io_in_valid_1(mesh_11_0_io_in_valid_1),
    .io_out_valid_0(mesh_11_0_io_out_valid_0),
    .io_out_valid_1(mesh_11_0_io_out_valid_1)
  );
  Tile mesh_11_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_1_clock),
    .io_in_a_0(mesh_11_1_io_in_a_0),
    .io_in_a_1(mesh_11_1_io_in_a_1),
    .io_in_b_0(mesh_11_1_io_in_b_0),
    .io_in_b_1(mesh_11_1_io_in_b_1),
    .io_in_d_0(mesh_11_1_io_in_d_0),
    .io_in_d_1(mesh_11_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_1_io_in_control_1_shift),
    .io_in_id_0(mesh_11_1_io_in_id_0),
    .io_in_id_1(mesh_11_1_io_in_id_1),
    .io_in_last_0(mesh_11_1_io_in_last_0),
    .io_in_last_1(mesh_11_1_io_in_last_1),
    .io_out_a_0(mesh_11_1_io_out_a_0),
    .io_out_a_1(mesh_11_1_io_out_a_1),
    .io_out_c_0(mesh_11_1_io_out_c_0),
    .io_out_c_1(mesh_11_1_io_out_c_1),
    .io_out_b_0(mesh_11_1_io_out_b_0),
    .io_out_b_1(mesh_11_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_1_io_out_control_1_shift),
    .io_out_id_0(mesh_11_1_io_out_id_0),
    .io_out_id_1(mesh_11_1_io_out_id_1),
    .io_out_last_0(mesh_11_1_io_out_last_0),
    .io_out_last_1(mesh_11_1_io_out_last_1),
    .io_in_valid_0(mesh_11_1_io_in_valid_0),
    .io_in_valid_1(mesh_11_1_io_in_valid_1),
    .io_out_valid_0(mesh_11_1_io_out_valid_0),
    .io_out_valid_1(mesh_11_1_io_out_valid_1)
  );
  Tile mesh_11_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_2_clock),
    .io_in_a_0(mesh_11_2_io_in_a_0),
    .io_in_a_1(mesh_11_2_io_in_a_1),
    .io_in_b_0(mesh_11_2_io_in_b_0),
    .io_in_b_1(mesh_11_2_io_in_b_1),
    .io_in_d_0(mesh_11_2_io_in_d_0),
    .io_in_d_1(mesh_11_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_2_io_in_control_1_shift),
    .io_in_id_0(mesh_11_2_io_in_id_0),
    .io_in_id_1(mesh_11_2_io_in_id_1),
    .io_in_last_0(mesh_11_2_io_in_last_0),
    .io_in_last_1(mesh_11_2_io_in_last_1),
    .io_out_a_0(mesh_11_2_io_out_a_0),
    .io_out_a_1(mesh_11_2_io_out_a_1),
    .io_out_c_0(mesh_11_2_io_out_c_0),
    .io_out_c_1(mesh_11_2_io_out_c_1),
    .io_out_b_0(mesh_11_2_io_out_b_0),
    .io_out_b_1(mesh_11_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_2_io_out_control_1_shift),
    .io_out_id_0(mesh_11_2_io_out_id_0),
    .io_out_id_1(mesh_11_2_io_out_id_1),
    .io_out_last_0(mesh_11_2_io_out_last_0),
    .io_out_last_1(mesh_11_2_io_out_last_1),
    .io_in_valid_0(mesh_11_2_io_in_valid_0),
    .io_in_valid_1(mesh_11_2_io_in_valid_1),
    .io_out_valid_0(mesh_11_2_io_out_valid_0),
    .io_out_valid_1(mesh_11_2_io_out_valid_1)
  );
  Tile mesh_11_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_3_clock),
    .io_in_a_0(mesh_11_3_io_in_a_0),
    .io_in_a_1(mesh_11_3_io_in_a_1),
    .io_in_b_0(mesh_11_3_io_in_b_0),
    .io_in_b_1(mesh_11_3_io_in_b_1),
    .io_in_d_0(mesh_11_3_io_in_d_0),
    .io_in_d_1(mesh_11_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_3_io_in_control_1_shift),
    .io_in_id_0(mesh_11_3_io_in_id_0),
    .io_in_id_1(mesh_11_3_io_in_id_1),
    .io_in_last_0(mesh_11_3_io_in_last_0),
    .io_in_last_1(mesh_11_3_io_in_last_1),
    .io_out_a_0(mesh_11_3_io_out_a_0),
    .io_out_a_1(mesh_11_3_io_out_a_1),
    .io_out_c_0(mesh_11_3_io_out_c_0),
    .io_out_c_1(mesh_11_3_io_out_c_1),
    .io_out_b_0(mesh_11_3_io_out_b_0),
    .io_out_b_1(mesh_11_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_3_io_out_control_1_shift),
    .io_out_id_0(mesh_11_3_io_out_id_0),
    .io_out_id_1(mesh_11_3_io_out_id_1),
    .io_out_last_0(mesh_11_3_io_out_last_0),
    .io_out_last_1(mesh_11_3_io_out_last_1),
    .io_in_valid_0(mesh_11_3_io_in_valid_0),
    .io_in_valid_1(mesh_11_3_io_in_valid_1),
    .io_out_valid_0(mesh_11_3_io_out_valid_0),
    .io_out_valid_1(mesh_11_3_io_out_valid_1)
  );
  Tile mesh_11_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_4_clock),
    .io_in_a_0(mesh_11_4_io_in_a_0),
    .io_in_a_1(mesh_11_4_io_in_a_1),
    .io_in_b_0(mesh_11_4_io_in_b_0),
    .io_in_b_1(mesh_11_4_io_in_b_1),
    .io_in_d_0(mesh_11_4_io_in_d_0),
    .io_in_d_1(mesh_11_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_4_io_in_control_1_shift),
    .io_in_id_0(mesh_11_4_io_in_id_0),
    .io_in_id_1(mesh_11_4_io_in_id_1),
    .io_in_last_0(mesh_11_4_io_in_last_0),
    .io_in_last_1(mesh_11_4_io_in_last_1),
    .io_out_a_0(mesh_11_4_io_out_a_0),
    .io_out_a_1(mesh_11_4_io_out_a_1),
    .io_out_c_0(mesh_11_4_io_out_c_0),
    .io_out_c_1(mesh_11_4_io_out_c_1),
    .io_out_b_0(mesh_11_4_io_out_b_0),
    .io_out_b_1(mesh_11_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_4_io_out_control_1_shift),
    .io_out_id_0(mesh_11_4_io_out_id_0),
    .io_out_id_1(mesh_11_4_io_out_id_1),
    .io_out_last_0(mesh_11_4_io_out_last_0),
    .io_out_last_1(mesh_11_4_io_out_last_1),
    .io_in_valid_0(mesh_11_4_io_in_valid_0),
    .io_in_valid_1(mesh_11_4_io_in_valid_1),
    .io_out_valid_0(mesh_11_4_io_out_valid_0),
    .io_out_valid_1(mesh_11_4_io_out_valid_1)
  );
  Tile mesh_11_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_5_clock),
    .io_in_a_0(mesh_11_5_io_in_a_0),
    .io_in_a_1(mesh_11_5_io_in_a_1),
    .io_in_b_0(mesh_11_5_io_in_b_0),
    .io_in_b_1(mesh_11_5_io_in_b_1),
    .io_in_d_0(mesh_11_5_io_in_d_0),
    .io_in_d_1(mesh_11_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_5_io_in_control_1_shift),
    .io_in_id_0(mesh_11_5_io_in_id_0),
    .io_in_id_1(mesh_11_5_io_in_id_1),
    .io_in_last_0(mesh_11_5_io_in_last_0),
    .io_in_last_1(mesh_11_5_io_in_last_1),
    .io_out_a_0(mesh_11_5_io_out_a_0),
    .io_out_a_1(mesh_11_5_io_out_a_1),
    .io_out_c_0(mesh_11_5_io_out_c_0),
    .io_out_c_1(mesh_11_5_io_out_c_1),
    .io_out_b_0(mesh_11_5_io_out_b_0),
    .io_out_b_1(mesh_11_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_5_io_out_control_1_shift),
    .io_out_id_0(mesh_11_5_io_out_id_0),
    .io_out_id_1(mesh_11_5_io_out_id_1),
    .io_out_last_0(mesh_11_5_io_out_last_0),
    .io_out_last_1(mesh_11_5_io_out_last_1),
    .io_in_valid_0(mesh_11_5_io_in_valid_0),
    .io_in_valid_1(mesh_11_5_io_in_valid_1),
    .io_out_valid_0(mesh_11_5_io_out_valid_0),
    .io_out_valid_1(mesh_11_5_io_out_valid_1)
  );
  Tile mesh_11_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_6_clock),
    .io_in_a_0(mesh_11_6_io_in_a_0),
    .io_in_a_1(mesh_11_6_io_in_a_1),
    .io_in_b_0(mesh_11_6_io_in_b_0),
    .io_in_b_1(mesh_11_6_io_in_b_1),
    .io_in_d_0(mesh_11_6_io_in_d_0),
    .io_in_d_1(mesh_11_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_6_io_in_control_1_shift),
    .io_in_id_0(mesh_11_6_io_in_id_0),
    .io_in_id_1(mesh_11_6_io_in_id_1),
    .io_in_last_0(mesh_11_6_io_in_last_0),
    .io_in_last_1(mesh_11_6_io_in_last_1),
    .io_out_a_0(mesh_11_6_io_out_a_0),
    .io_out_a_1(mesh_11_6_io_out_a_1),
    .io_out_c_0(mesh_11_6_io_out_c_0),
    .io_out_c_1(mesh_11_6_io_out_c_1),
    .io_out_b_0(mesh_11_6_io_out_b_0),
    .io_out_b_1(mesh_11_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_6_io_out_control_1_shift),
    .io_out_id_0(mesh_11_6_io_out_id_0),
    .io_out_id_1(mesh_11_6_io_out_id_1),
    .io_out_last_0(mesh_11_6_io_out_last_0),
    .io_out_last_1(mesh_11_6_io_out_last_1),
    .io_in_valid_0(mesh_11_6_io_in_valid_0),
    .io_in_valid_1(mesh_11_6_io_in_valid_1),
    .io_out_valid_0(mesh_11_6_io_out_valid_0),
    .io_out_valid_1(mesh_11_6_io_out_valid_1)
  );
  Tile mesh_11_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_7_clock),
    .io_in_a_0(mesh_11_7_io_in_a_0),
    .io_in_a_1(mesh_11_7_io_in_a_1),
    .io_in_b_0(mesh_11_7_io_in_b_0),
    .io_in_b_1(mesh_11_7_io_in_b_1),
    .io_in_d_0(mesh_11_7_io_in_d_0),
    .io_in_d_1(mesh_11_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_7_io_in_control_1_shift),
    .io_in_id_0(mesh_11_7_io_in_id_0),
    .io_in_id_1(mesh_11_7_io_in_id_1),
    .io_in_last_0(mesh_11_7_io_in_last_0),
    .io_in_last_1(mesh_11_7_io_in_last_1),
    .io_out_a_0(mesh_11_7_io_out_a_0),
    .io_out_a_1(mesh_11_7_io_out_a_1),
    .io_out_c_0(mesh_11_7_io_out_c_0),
    .io_out_c_1(mesh_11_7_io_out_c_1),
    .io_out_b_0(mesh_11_7_io_out_b_0),
    .io_out_b_1(mesh_11_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_7_io_out_control_1_shift),
    .io_out_id_0(mesh_11_7_io_out_id_0),
    .io_out_id_1(mesh_11_7_io_out_id_1),
    .io_out_last_0(mesh_11_7_io_out_last_0),
    .io_out_last_1(mesh_11_7_io_out_last_1),
    .io_in_valid_0(mesh_11_7_io_in_valid_0),
    .io_in_valid_1(mesh_11_7_io_in_valid_1),
    .io_out_valid_0(mesh_11_7_io_out_valid_0),
    .io_out_valid_1(mesh_11_7_io_out_valid_1)
  );
  Tile mesh_11_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_8_clock),
    .io_in_a_0(mesh_11_8_io_in_a_0),
    .io_in_a_1(mesh_11_8_io_in_a_1),
    .io_in_b_0(mesh_11_8_io_in_b_0),
    .io_in_b_1(mesh_11_8_io_in_b_1),
    .io_in_d_0(mesh_11_8_io_in_d_0),
    .io_in_d_1(mesh_11_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_8_io_in_control_1_shift),
    .io_in_id_0(mesh_11_8_io_in_id_0),
    .io_in_id_1(mesh_11_8_io_in_id_1),
    .io_in_last_0(mesh_11_8_io_in_last_0),
    .io_in_last_1(mesh_11_8_io_in_last_1),
    .io_out_a_0(mesh_11_8_io_out_a_0),
    .io_out_a_1(mesh_11_8_io_out_a_1),
    .io_out_c_0(mesh_11_8_io_out_c_0),
    .io_out_c_1(mesh_11_8_io_out_c_1),
    .io_out_b_0(mesh_11_8_io_out_b_0),
    .io_out_b_1(mesh_11_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_8_io_out_control_1_shift),
    .io_out_id_0(mesh_11_8_io_out_id_0),
    .io_out_id_1(mesh_11_8_io_out_id_1),
    .io_out_last_0(mesh_11_8_io_out_last_0),
    .io_out_last_1(mesh_11_8_io_out_last_1),
    .io_in_valid_0(mesh_11_8_io_in_valid_0),
    .io_in_valid_1(mesh_11_8_io_in_valid_1),
    .io_out_valid_0(mesh_11_8_io_out_valid_0),
    .io_out_valid_1(mesh_11_8_io_out_valid_1)
  );
  Tile mesh_11_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_9_clock),
    .io_in_a_0(mesh_11_9_io_in_a_0),
    .io_in_a_1(mesh_11_9_io_in_a_1),
    .io_in_b_0(mesh_11_9_io_in_b_0),
    .io_in_b_1(mesh_11_9_io_in_b_1),
    .io_in_d_0(mesh_11_9_io_in_d_0),
    .io_in_d_1(mesh_11_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_9_io_in_control_1_shift),
    .io_in_id_0(mesh_11_9_io_in_id_0),
    .io_in_id_1(mesh_11_9_io_in_id_1),
    .io_in_last_0(mesh_11_9_io_in_last_0),
    .io_in_last_1(mesh_11_9_io_in_last_1),
    .io_out_a_0(mesh_11_9_io_out_a_0),
    .io_out_a_1(mesh_11_9_io_out_a_1),
    .io_out_c_0(mesh_11_9_io_out_c_0),
    .io_out_c_1(mesh_11_9_io_out_c_1),
    .io_out_b_0(mesh_11_9_io_out_b_0),
    .io_out_b_1(mesh_11_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_9_io_out_control_1_shift),
    .io_out_id_0(mesh_11_9_io_out_id_0),
    .io_out_id_1(mesh_11_9_io_out_id_1),
    .io_out_last_0(mesh_11_9_io_out_last_0),
    .io_out_last_1(mesh_11_9_io_out_last_1),
    .io_in_valid_0(mesh_11_9_io_in_valid_0),
    .io_in_valid_1(mesh_11_9_io_in_valid_1),
    .io_out_valid_0(mesh_11_9_io_out_valid_0),
    .io_out_valid_1(mesh_11_9_io_out_valid_1)
  );
  Tile mesh_11_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_10_clock),
    .io_in_a_0(mesh_11_10_io_in_a_0),
    .io_in_a_1(mesh_11_10_io_in_a_1),
    .io_in_b_0(mesh_11_10_io_in_b_0),
    .io_in_b_1(mesh_11_10_io_in_b_1),
    .io_in_d_0(mesh_11_10_io_in_d_0),
    .io_in_d_1(mesh_11_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_10_io_in_control_1_shift),
    .io_in_id_0(mesh_11_10_io_in_id_0),
    .io_in_id_1(mesh_11_10_io_in_id_1),
    .io_in_last_0(mesh_11_10_io_in_last_0),
    .io_in_last_1(mesh_11_10_io_in_last_1),
    .io_out_a_0(mesh_11_10_io_out_a_0),
    .io_out_a_1(mesh_11_10_io_out_a_1),
    .io_out_c_0(mesh_11_10_io_out_c_0),
    .io_out_c_1(mesh_11_10_io_out_c_1),
    .io_out_b_0(mesh_11_10_io_out_b_0),
    .io_out_b_1(mesh_11_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_10_io_out_control_1_shift),
    .io_out_id_0(mesh_11_10_io_out_id_0),
    .io_out_id_1(mesh_11_10_io_out_id_1),
    .io_out_last_0(mesh_11_10_io_out_last_0),
    .io_out_last_1(mesh_11_10_io_out_last_1),
    .io_in_valid_0(mesh_11_10_io_in_valid_0),
    .io_in_valid_1(mesh_11_10_io_in_valid_1),
    .io_out_valid_0(mesh_11_10_io_out_valid_0),
    .io_out_valid_1(mesh_11_10_io_out_valid_1)
  );
  Tile mesh_11_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_11_clock),
    .io_in_a_0(mesh_11_11_io_in_a_0),
    .io_in_a_1(mesh_11_11_io_in_a_1),
    .io_in_b_0(mesh_11_11_io_in_b_0),
    .io_in_b_1(mesh_11_11_io_in_b_1),
    .io_in_d_0(mesh_11_11_io_in_d_0),
    .io_in_d_1(mesh_11_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_11_io_in_control_1_shift),
    .io_in_id_0(mesh_11_11_io_in_id_0),
    .io_in_id_1(mesh_11_11_io_in_id_1),
    .io_in_last_0(mesh_11_11_io_in_last_0),
    .io_in_last_1(mesh_11_11_io_in_last_1),
    .io_out_a_0(mesh_11_11_io_out_a_0),
    .io_out_a_1(mesh_11_11_io_out_a_1),
    .io_out_c_0(mesh_11_11_io_out_c_0),
    .io_out_c_1(mesh_11_11_io_out_c_1),
    .io_out_b_0(mesh_11_11_io_out_b_0),
    .io_out_b_1(mesh_11_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_11_io_out_control_1_shift),
    .io_out_id_0(mesh_11_11_io_out_id_0),
    .io_out_id_1(mesh_11_11_io_out_id_1),
    .io_out_last_0(mesh_11_11_io_out_last_0),
    .io_out_last_1(mesh_11_11_io_out_last_1),
    .io_in_valid_0(mesh_11_11_io_in_valid_0),
    .io_in_valid_1(mesh_11_11_io_in_valid_1),
    .io_out_valid_0(mesh_11_11_io_out_valid_0),
    .io_out_valid_1(mesh_11_11_io_out_valid_1)
  );
  Tile mesh_11_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_12_clock),
    .io_in_a_0(mesh_11_12_io_in_a_0),
    .io_in_a_1(mesh_11_12_io_in_a_1),
    .io_in_b_0(mesh_11_12_io_in_b_0),
    .io_in_b_1(mesh_11_12_io_in_b_1),
    .io_in_d_0(mesh_11_12_io_in_d_0),
    .io_in_d_1(mesh_11_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_12_io_in_control_1_shift),
    .io_in_id_0(mesh_11_12_io_in_id_0),
    .io_in_id_1(mesh_11_12_io_in_id_1),
    .io_in_last_0(mesh_11_12_io_in_last_0),
    .io_in_last_1(mesh_11_12_io_in_last_1),
    .io_out_a_0(mesh_11_12_io_out_a_0),
    .io_out_a_1(mesh_11_12_io_out_a_1),
    .io_out_c_0(mesh_11_12_io_out_c_0),
    .io_out_c_1(mesh_11_12_io_out_c_1),
    .io_out_b_0(mesh_11_12_io_out_b_0),
    .io_out_b_1(mesh_11_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_12_io_out_control_1_shift),
    .io_out_id_0(mesh_11_12_io_out_id_0),
    .io_out_id_1(mesh_11_12_io_out_id_1),
    .io_out_last_0(mesh_11_12_io_out_last_0),
    .io_out_last_1(mesh_11_12_io_out_last_1),
    .io_in_valid_0(mesh_11_12_io_in_valid_0),
    .io_in_valid_1(mesh_11_12_io_in_valid_1),
    .io_out_valid_0(mesh_11_12_io_out_valid_0),
    .io_out_valid_1(mesh_11_12_io_out_valid_1)
  );
  Tile mesh_11_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_13_clock),
    .io_in_a_0(mesh_11_13_io_in_a_0),
    .io_in_a_1(mesh_11_13_io_in_a_1),
    .io_in_b_0(mesh_11_13_io_in_b_0),
    .io_in_b_1(mesh_11_13_io_in_b_1),
    .io_in_d_0(mesh_11_13_io_in_d_0),
    .io_in_d_1(mesh_11_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_13_io_in_control_1_shift),
    .io_in_id_0(mesh_11_13_io_in_id_0),
    .io_in_id_1(mesh_11_13_io_in_id_1),
    .io_in_last_0(mesh_11_13_io_in_last_0),
    .io_in_last_1(mesh_11_13_io_in_last_1),
    .io_out_a_0(mesh_11_13_io_out_a_0),
    .io_out_a_1(mesh_11_13_io_out_a_1),
    .io_out_c_0(mesh_11_13_io_out_c_0),
    .io_out_c_1(mesh_11_13_io_out_c_1),
    .io_out_b_0(mesh_11_13_io_out_b_0),
    .io_out_b_1(mesh_11_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_13_io_out_control_1_shift),
    .io_out_id_0(mesh_11_13_io_out_id_0),
    .io_out_id_1(mesh_11_13_io_out_id_1),
    .io_out_last_0(mesh_11_13_io_out_last_0),
    .io_out_last_1(mesh_11_13_io_out_last_1),
    .io_in_valid_0(mesh_11_13_io_in_valid_0),
    .io_in_valid_1(mesh_11_13_io_in_valid_1),
    .io_out_valid_0(mesh_11_13_io_out_valid_0),
    .io_out_valid_1(mesh_11_13_io_out_valid_1)
  );
  Tile mesh_11_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_14_clock),
    .io_in_a_0(mesh_11_14_io_in_a_0),
    .io_in_a_1(mesh_11_14_io_in_a_1),
    .io_in_b_0(mesh_11_14_io_in_b_0),
    .io_in_b_1(mesh_11_14_io_in_b_1),
    .io_in_d_0(mesh_11_14_io_in_d_0),
    .io_in_d_1(mesh_11_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_14_io_in_control_1_shift),
    .io_in_id_0(mesh_11_14_io_in_id_0),
    .io_in_id_1(mesh_11_14_io_in_id_1),
    .io_in_last_0(mesh_11_14_io_in_last_0),
    .io_in_last_1(mesh_11_14_io_in_last_1),
    .io_out_a_0(mesh_11_14_io_out_a_0),
    .io_out_a_1(mesh_11_14_io_out_a_1),
    .io_out_c_0(mesh_11_14_io_out_c_0),
    .io_out_c_1(mesh_11_14_io_out_c_1),
    .io_out_b_0(mesh_11_14_io_out_b_0),
    .io_out_b_1(mesh_11_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_14_io_out_control_1_shift),
    .io_out_id_0(mesh_11_14_io_out_id_0),
    .io_out_id_1(mesh_11_14_io_out_id_1),
    .io_out_last_0(mesh_11_14_io_out_last_0),
    .io_out_last_1(mesh_11_14_io_out_last_1),
    .io_in_valid_0(mesh_11_14_io_in_valid_0),
    .io_in_valid_1(mesh_11_14_io_in_valid_1),
    .io_out_valid_0(mesh_11_14_io_out_valid_0),
    .io_out_valid_1(mesh_11_14_io_out_valid_1)
  );
  Tile mesh_11_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_11_15_clock),
    .io_in_a_0(mesh_11_15_io_in_a_0),
    .io_in_a_1(mesh_11_15_io_in_a_1),
    .io_in_b_0(mesh_11_15_io_in_b_0),
    .io_in_b_1(mesh_11_15_io_in_b_1),
    .io_in_d_0(mesh_11_15_io_in_d_0),
    .io_in_d_1(mesh_11_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_11_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_11_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_11_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_11_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_11_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_11_15_io_in_control_1_shift),
    .io_in_id_0(mesh_11_15_io_in_id_0),
    .io_in_id_1(mesh_11_15_io_in_id_1),
    .io_in_last_0(mesh_11_15_io_in_last_0),
    .io_in_last_1(mesh_11_15_io_in_last_1),
    .io_out_a_0(mesh_11_15_io_out_a_0),
    .io_out_a_1(mesh_11_15_io_out_a_1),
    .io_out_c_0(mesh_11_15_io_out_c_0),
    .io_out_c_1(mesh_11_15_io_out_c_1),
    .io_out_b_0(mesh_11_15_io_out_b_0),
    .io_out_b_1(mesh_11_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_11_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_11_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_11_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_11_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_11_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_11_15_io_out_control_1_shift),
    .io_out_id_0(mesh_11_15_io_out_id_0),
    .io_out_id_1(mesh_11_15_io_out_id_1),
    .io_out_last_0(mesh_11_15_io_out_last_0),
    .io_out_last_1(mesh_11_15_io_out_last_1),
    .io_in_valid_0(mesh_11_15_io_in_valid_0),
    .io_in_valid_1(mesh_11_15_io_in_valid_1),
    .io_out_valid_0(mesh_11_15_io_out_valid_0),
    .io_out_valid_1(mesh_11_15_io_out_valid_1)
  );
  Tile mesh_12_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_0_clock),
    .io_in_a_0(mesh_12_0_io_in_a_0),
    .io_in_a_1(mesh_12_0_io_in_a_1),
    .io_in_b_0(mesh_12_0_io_in_b_0),
    .io_in_b_1(mesh_12_0_io_in_b_1),
    .io_in_d_0(mesh_12_0_io_in_d_0),
    .io_in_d_1(mesh_12_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_0_io_in_control_1_shift),
    .io_in_id_0(mesh_12_0_io_in_id_0),
    .io_in_id_1(mesh_12_0_io_in_id_1),
    .io_in_last_0(mesh_12_0_io_in_last_0),
    .io_in_last_1(mesh_12_0_io_in_last_1),
    .io_out_a_0(mesh_12_0_io_out_a_0),
    .io_out_a_1(mesh_12_0_io_out_a_1),
    .io_out_c_0(mesh_12_0_io_out_c_0),
    .io_out_c_1(mesh_12_0_io_out_c_1),
    .io_out_b_0(mesh_12_0_io_out_b_0),
    .io_out_b_1(mesh_12_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_0_io_out_control_1_shift),
    .io_out_id_0(mesh_12_0_io_out_id_0),
    .io_out_id_1(mesh_12_0_io_out_id_1),
    .io_out_last_0(mesh_12_0_io_out_last_0),
    .io_out_last_1(mesh_12_0_io_out_last_1),
    .io_in_valid_0(mesh_12_0_io_in_valid_0),
    .io_in_valid_1(mesh_12_0_io_in_valid_1),
    .io_out_valid_0(mesh_12_0_io_out_valid_0),
    .io_out_valid_1(mesh_12_0_io_out_valid_1)
  );
  Tile mesh_12_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_1_clock),
    .io_in_a_0(mesh_12_1_io_in_a_0),
    .io_in_a_1(mesh_12_1_io_in_a_1),
    .io_in_b_0(mesh_12_1_io_in_b_0),
    .io_in_b_1(mesh_12_1_io_in_b_1),
    .io_in_d_0(mesh_12_1_io_in_d_0),
    .io_in_d_1(mesh_12_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_1_io_in_control_1_shift),
    .io_in_id_0(mesh_12_1_io_in_id_0),
    .io_in_id_1(mesh_12_1_io_in_id_1),
    .io_in_last_0(mesh_12_1_io_in_last_0),
    .io_in_last_1(mesh_12_1_io_in_last_1),
    .io_out_a_0(mesh_12_1_io_out_a_0),
    .io_out_a_1(mesh_12_1_io_out_a_1),
    .io_out_c_0(mesh_12_1_io_out_c_0),
    .io_out_c_1(mesh_12_1_io_out_c_1),
    .io_out_b_0(mesh_12_1_io_out_b_0),
    .io_out_b_1(mesh_12_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_1_io_out_control_1_shift),
    .io_out_id_0(mesh_12_1_io_out_id_0),
    .io_out_id_1(mesh_12_1_io_out_id_1),
    .io_out_last_0(mesh_12_1_io_out_last_0),
    .io_out_last_1(mesh_12_1_io_out_last_1),
    .io_in_valid_0(mesh_12_1_io_in_valid_0),
    .io_in_valid_1(mesh_12_1_io_in_valid_1),
    .io_out_valid_0(mesh_12_1_io_out_valid_0),
    .io_out_valid_1(mesh_12_1_io_out_valid_1)
  );
  Tile mesh_12_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_2_clock),
    .io_in_a_0(mesh_12_2_io_in_a_0),
    .io_in_a_1(mesh_12_2_io_in_a_1),
    .io_in_b_0(mesh_12_2_io_in_b_0),
    .io_in_b_1(mesh_12_2_io_in_b_1),
    .io_in_d_0(mesh_12_2_io_in_d_0),
    .io_in_d_1(mesh_12_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_2_io_in_control_1_shift),
    .io_in_id_0(mesh_12_2_io_in_id_0),
    .io_in_id_1(mesh_12_2_io_in_id_1),
    .io_in_last_0(mesh_12_2_io_in_last_0),
    .io_in_last_1(mesh_12_2_io_in_last_1),
    .io_out_a_0(mesh_12_2_io_out_a_0),
    .io_out_a_1(mesh_12_2_io_out_a_1),
    .io_out_c_0(mesh_12_2_io_out_c_0),
    .io_out_c_1(mesh_12_2_io_out_c_1),
    .io_out_b_0(mesh_12_2_io_out_b_0),
    .io_out_b_1(mesh_12_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_2_io_out_control_1_shift),
    .io_out_id_0(mesh_12_2_io_out_id_0),
    .io_out_id_1(mesh_12_2_io_out_id_1),
    .io_out_last_0(mesh_12_2_io_out_last_0),
    .io_out_last_1(mesh_12_2_io_out_last_1),
    .io_in_valid_0(mesh_12_2_io_in_valid_0),
    .io_in_valid_1(mesh_12_2_io_in_valid_1),
    .io_out_valid_0(mesh_12_2_io_out_valid_0),
    .io_out_valid_1(mesh_12_2_io_out_valid_1)
  );
  Tile mesh_12_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_3_clock),
    .io_in_a_0(mesh_12_3_io_in_a_0),
    .io_in_a_1(mesh_12_3_io_in_a_1),
    .io_in_b_0(mesh_12_3_io_in_b_0),
    .io_in_b_1(mesh_12_3_io_in_b_1),
    .io_in_d_0(mesh_12_3_io_in_d_0),
    .io_in_d_1(mesh_12_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_3_io_in_control_1_shift),
    .io_in_id_0(mesh_12_3_io_in_id_0),
    .io_in_id_1(mesh_12_3_io_in_id_1),
    .io_in_last_0(mesh_12_3_io_in_last_0),
    .io_in_last_1(mesh_12_3_io_in_last_1),
    .io_out_a_0(mesh_12_3_io_out_a_0),
    .io_out_a_1(mesh_12_3_io_out_a_1),
    .io_out_c_0(mesh_12_3_io_out_c_0),
    .io_out_c_1(mesh_12_3_io_out_c_1),
    .io_out_b_0(mesh_12_3_io_out_b_0),
    .io_out_b_1(mesh_12_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_3_io_out_control_1_shift),
    .io_out_id_0(mesh_12_3_io_out_id_0),
    .io_out_id_1(mesh_12_3_io_out_id_1),
    .io_out_last_0(mesh_12_3_io_out_last_0),
    .io_out_last_1(mesh_12_3_io_out_last_1),
    .io_in_valid_0(mesh_12_3_io_in_valid_0),
    .io_in_valid_1(mesh_12_3_io_in_valid_1),
    .io_out_valid_0(mesh_12_3_io_out_valid_0),
    .io_out_valid_1(mesh_12_3_io_out_valid_1)
  );
  Tile mesh_12_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_4_clock),
    .io_in_a_0(mesh_12_4_io_in_a_0),
    .io_in_a_1(mesh_12_4_io_in_a_1),
    .io_in_b_0(mesh_12_4_io_in_b_0),
    .io_in_b_1(mesh_12_4_io_in_b_1),
    .io_in_d_0(mesh_12_4_io_in_d_0),
    .io_in_d_1(mesh_12_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_4_io_in_control_1_shift),
    .io_in_id_0(mesh_12_4_io_in_id_0),
    .io_in_id_1(mesh_12_4_io_in_id_1),
    .io_in_last_0(mesh_12_4_io_in_last_0),
    .io_in_last_1(mesh_12_4_io_in_last_1),
    .io_out_a_0(mesh_12_4_io_out_a_0),
    .io_out_a_1(mesh_12_4_io_out_a_1),
    .io_out_c_0(mesh_12_4_io_out_c_0),
    .io_out_c_1(mesh_12_4_io_out_c_1),
    .io_out_b_0(mesh_12_4_io_out_b_0),
    .io_out_b_1(mesh_12_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_4_io_out_control_1_shift),
    .io_out_id_0(mesh_12_4_io_out_id_0),
    .io_out_id_1(mesh_12_4_io_out_id_1),
    .io_out_last_0(mesh_12_4_io_out_last_0),
    .io_out_last_1(mesh_12_4_io_out_last_1),
    .io_in_valid_0(mesh_12_4_io_in_valid_0),
    .io_in_valid_1(mesh_12_4_io_in_valid_1),
    .io_out_valid_0(mesh_12_4_io_out_valid_0),
    .io_out_valid_1(mesh_12_4_io_out_valid_1)
  );
  Tile mesh_12_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_5_clock),
    .io_in_a_0(mesh_12_5_io_in_a_0),
    .io_in_a_1(mesh_12_5_io_in_a_1),
    .io_in_b_0(mesh_12_5_io_in_b_0),
    .io_in_b_1(mesh_12_5_io_in_b_1),
    .io_in_d_0(mesh_12_5_io_in_d_0),
    .io_in_d_1(mesh_12_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_5_io_in_control_1_shift),
    .io_in_id_0(mesh_12_5_io_in_id_0),
    .io_in_id_1(mesh_12_5_io_in_id_1),
    .io_in_last_0(mesh_12_5_io_in_last_0),
    .io_in_last_1(mesh_12_5_io_in_last_1),
    .io_out_a_0(mesh_12_5_io_out_a_0),
    .io_out_a_1(mesh_12_5_io_out_a_1),
    .io_out_c_0(mesh_12_5_io_out_c_0),
    .io_out_c_1(mesh_12_5_io_out_c_1),
    .io_out_b_0(mesh_12_5_io_out_b_0),
    .io_out_b_1(mesh_12_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_5_io_out_control_1_shift),
    .io_out_id_0(mesh_12_5_io_out_id_0),
    .io_out_id_1(mesh_12_5_io_out_id_1),
    .io_out_last_0(mesh_12_5_io_out_last_0),
    .io_out_last_1(mesh_12_5_io_out_last_1),
    .io_in_valid_0(mesh_12_5_io_in_valid_0),
    .io_in_valid_1(mesh_12_5_io_in_valid_1),
    .io_out_valid_0(mesh_12_5_io_out_valid_0),
    .io_out_valid_1(mesh_12_5_io_out_valid_1)
  );
  Tile mesh_12_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_6_clock),
    .io_in_a_0(mesh_12_6_io_in_a_0),
    .io_in_a_1(mesh_12_6_io_in_a_1),
    .io_in_b_0(mesh_12_6_io_in_b_0),
    .io_in_b_1(mesh_12_6_io_in_b_1),
    .io_in_d_0(mesh_12_6_io_in_d_0),
    .io_in_d_1(mesh_12_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_6_io_in_control_1_shift),
    .io_in_id_0(mesh_12_6_io_in_id_0),
    .io_in_id_1(mesh_12_6_io_in_id_1),
    .io_in_last_0(mesh_12_6_io_in_last_0),
    .io_in_last_1(mesh_12_6_io_in_last_1),
    .io_out_a_0(mesh_12_6_io_out_a_0),
    .io_out_a_1(mesh_12_6_io_out_a_1),
    .io_out_c_0(mesh_12_6_io_out_c_0),
    .io_out_c_1(mesh_12_6_io_out_c_1),
    .io_out_b_0(mesh_12_6_io_out_b_0),
    .io_out_b_1(mesh_12_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_6_io_out_control_1_shift),
    .io_out_id_0(mesh_12_6_io_out_id_0),
    .io_out_id_1(mesh_12_6_io_out_id_1),
    .io_out_last_0(mesh_12_6_io_out_last_0),
    .io_out_last_1(mesh_12_6_io_out_last_1),
    .io_in_valid_0(mesh_12_6_io_in_valid_0),
    .io_in_valid_1(mesh_12_6_io_in_valid_1),
    .io_out_valid_0(mesh_12_6_io_out_valid_0),
    .io_out_valid_1(mesh_12_6_io_out_valid_1)
  );
  Tile mesh_12_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_7_clock),
    .io_in_a_0(mesh_12_7_io_in_a_0),
    .io_in_a_1(mesh_12_7_io_in_a_1),
    .io_in_b_0(mesh_12_7_io_in_b_0),
    .io_in_b_1(mesh_12_7_io_in_b_1),
    .io_in_d_0(mesh_12_7_io_in_d_0),
    .io_in_d_1(mesh_12_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_7_io_in_control_1_shift),
    .io_in_id_0(mesh_12_7_io_in_id_0),
    .io_in_id_1(mesh_12_7_io_in_id_1),
    .io_in_last_0(mesh_12_7_io_in_last_0),
    .io_in_last_1(mesh_12_7_io_in_last_1),
    .io_out_a_0(mesh_12_7_io_out_a_0),
    .io_out_a_1(mesh_12_7_io_out_a_1),
    .io_out_c_0(mesh_12_7_io_out_c_0),
    .io_out_c_1(mesh_12_7_io_out_c_1),
    .io_out_b_0(mesh_12_7_io_out_b_0),
    .io_out_b_1(mesh_12_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_7_io_out_control_1_shift),
    .io_out_id_0(mesh_12_7_io_out_id_0),
    .io_out_id_1(mesh_12_7_io_out_id_1),
    .io_out_last_0(mesh_12_7_io_out_last_0),
    .io_out_last_1(mesh_12_7_io_out_last_1),
    .io_in_valid_0(mesh_12_7_io_in_valid_0),
    .io_in_valid_1(mesh_12_7_io_in_valid_1),
    .io_out_valid_0(mesh_12_7_io_out_valid_0),
    .io_out_valid_1(mesh_12_7_io_out_valid_1)
  );
  Tile mesh_12_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_8_clock),
    .io_in_a_0(mesh_12_8_io_in_a_0),
    .io_in_a_1(mesh_12_8_io_in_a_1),
    .io_in_b_0(mesh_12_8_io_in_b_0),
    .io_in_b_1(mesh_12_8_io_in_b_1),
    .io_in_d_0(mesh_12_8_io_in_d_0),
    .io_in_d_1(mesh_12_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_8_io_in_control_1_shift),
    .io_in_id_0(mesh_12_8_io_in_id_0),
    .io_in_id_1(mesh_12_8_io_in_id_1),
    .io_in_last_0(mesh_12_8_io_in_last_0),
    .io_in_last_1(mesh_12_8_io_in_last_1),
    .io_out_a_0(mesh_12_8_io_out_a_0),
    .io_out_a_1(mesh_12_8_io_out_a_1),
    .io_out_c_0(mesh_12_8_io_out_c_0),
    .io_out_c_1(mesh_12_8_io_out_c_1),
    .io_out_b_0(mesh_12_8_io_out_b_0),
    .io_out_b_1(mesh_12_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_8_io_out_control_1_shift),
    .io_out_id_0(mesh_12_8_io_out_id_0),
    .io_out_id_1(mesh_12_8_io_out_id_1),
    .io_out_last_0(mesh_12_8_io_out_last_0),
    .io_out_last_1(mesh_12_8_io_out_last_1),
    .io_in_valid_0(mesh_12_8_io_in_valid_0),
    .io_in_valid_1(mesh_12_8_io_in_valid_1),
    .io_out_valid_0(mesh_12_8_io_out_valid_0),
    .io_out_valid_1(mesh_12_8_io_out_valid_1)
  );
  Tile mesh_12_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_9_clock),
    .io_in_a_0(mesh_12_9_io_in_a_0),
    .io_in_a_1(mesh_12_9_io_in_a_1),
    .io_in_b_0(mesh_12_9_io_in_b_0),
    .io_in_b_1(mesh_12_9_io_in_b_1),
    .io_in_d_0(mesh_12_9_io_in_d_0),
    .io_in_d_1(mesh_12_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_9_io_in_control_1_shift),
    .io_in_id_0(mesh_12_9_io_in_id_0),
    .io_in_id_1(mesh_12_9_io_in_id_1),
    .io_in_last_0(mesh_12_9_io_in_last_0),
    .io_in_last_1(mesh_12_9_io_in_last_1),
    .io_out_a_0(mesh_12_9_io_out_a_0),
    .io_out_a_1(mesh_12_9_io_out_a_1),
    .io_out_c_0(mesh_12_9_io_out_c_0),
    .io_out_c_1(mesh_12_9_io_out_c_1),
    .io_out_b_0(mesh_12_9_io_out_b_0),
    .io_out_b_1(mesh_12_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_9_io_out_control_1_shift),
    .io_out_id_0(mesh_12_9_io_out_id_0),
    .io_out_id_1(mesh_12_9_io_out_id_1),
    .io_out_last_0(mesh_12_9_io_out_last_0),
    .io_out_last_1(mesh_12_9_io_out_last_1),
    .io_in_valid_0(mesh_12_9_io_in_valid_0),
    .io_in_valid_1(mesh_12_9_io_in_valid_1),
    .io_out_valid_0(mesh_12_9_io_out_valid_0),
    .io_out_valid_1(mesh_12_9_io_out_valid_1)
  );
  Tile mesh_12_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_10_clock),
    .io_in_a_0(mesh_12_10_io_in_a_0),
    .io_in_a_1(mesh_12_10_io_in_a_1),
    .io_in_b_0(mesh_12_10_io_in_b_0),
    .io_in_b_1(mesh_12_10_io_in_b_1),
    .io_in_d_0(mesh_12_10_io_in_d_0),
    .io_in_d_1(mesh_12_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_10_io_in_control_1_shift),
    .io_in_id_0(mesh_12_10_io_in_id_0),
    .io_in_id_1(mesh_12_10_io_in_id_1),
    .io_in_last_0(mesh_12_10_io_in_last_0),
    .io_in_last_1(mesh_12_10_io_in_last_1),
    .io_out_a_0(mesh_12_10_io_out_a_0),
    .io_out_a_1(mesh_12_10_io_out_a_1),
    .io_out_c_0(mesh_12_10_io_out_c_0),
    .io_out_c_1(mesh_12_10_io_out_c_1),
    .io_out_b_0(mesh_12_10_io_out_b_0),
    .io_out_b_1(mesh_12_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_10_io_out_control_1_shift),
    .io_out_id_0(mesh_12_10_io_out_id_0),
    .io_out_id_1(mesh_12_10_io_out_id_1),
    .io_out_last_0(mesh_12_10_io_out_last_0),
    .io_out_last_1(mesh_12_10_io_out_last_1),
    .io_in_valid_0(mesh_12_10_io_in_valid_0),
    .io_in_valid_1(mesh_12_10_io_in_valid_1),
    .io_out_valid_0(mesh_12_10_io_out_valid_0),
    .io_out_valid_1(mesh_12_10_io_out_valid_1)
  );
  Tile mesh_12_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_11_clock),
    .io_in_a_0(mesh_12_11_io_in_a_0),
    .io_in_a_1(mesh_12_11_io_in_a_1),
    .io_in_b_0(mesh_12_11_io_in_b_0),
    .io_in_b_1(mesh_12_11_io_in_b_1),
    .io_in_d_0(mesh_12_11_io_in_d_0),
    .io_in_d_1(mesh_12_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_11_io_in_control_1_shift),
    .io_in_id_0(mesh_12_11_io_in_id_0),
    .io_in_id_1(mesh_12_11_io_in_id_1),
    .io_in_last_0(mesh_12_11_io_in_last_0),
    .io_in_last_1(mesh_12_11_io_in_last_1),
    .io_out_a_0(mesh_12_11_io_out_a_0),
    .io_out_a_1(mesh_12_11_io_out_a_1),
    .io_out_c_0(mesh_12_11_io_out_c_0),
    .io_out_c_1(mesh_12_11_io_out_c_1),
    .io_out_b_0(mesh_12_11_io_out_b_0),
    .io_out_b_1(mesh_12_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_11_io_out_control_1_shift),
    .io_out_id_0(mesh_12_11_io_out_id_0),
    .io_out_id_1(mesh_12_11_io_out_id_1),
    .io_out_last_0(mesh_12_11_io_out_last_0),
    .io_out_last_1(mesh_12_11_io_out_last_1),
    .io_in_valid_0(mesh_12_11_io_in_valid_0),
    .io_in_valid_1(mesh_12_11_io_in_valid_1),
    .io_out_valid_0(mesh_12_11_io_out_valid_0),
    .io_out_valid_1(mesh_12_11_io_out_valid_1)
  );
  Tile mesh_12_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_12_clock),
    .io_in_a_0(mesh_12_12_io_in_a_0),
    .io_in_a_1(mesh_12_12_io_in_a_1),
    .io_in_b_0(mesh_12_12_io_in_b_0),
    .io_in_b_1(mesh_12_12_io_in_b_1),
    .io_in_d_0(mesh_12_12_io_in_d_0),
    .io_in_d_1(mesh_12_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_12_io_in_control_1_shift),
    .io_in_id_0(mesh_12_12_io_in_id_0),
    .io_in_id_1(mesh_12_12_io_in_id_1),
    .io_in_last_0(mesh_12_12_io_in_last_0),
    .io_in_last_1(mesh_12_12_io_in_last_1),
    .io_out_a_0(mesh_12_12_io_out_a_0),
    .io_out_a_1(mesh_12_12_io_out_a_1),
    .io_out_c_0(mesh_12_12_io_out_c_0),
    .io_out_c_1(mesh_12_12_io_out_c_1),
    .io_out_b_0(mesh_12_12_io_out_b_0),
    .io_out_b_1(mesh_12_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_12_io_out_control_1_shift),
    .io_out_id_0(mesh_12_12_io_out_id_0),
    .io_out_id_1(mesh_12_12_io_out_id_1),
    .io_out_last_0(mesh_12_12_io_out_last_0),
    .io_out_last_1(mesh_12_12_io_out_last_1),
    .io_in_valid_0(mesh_12_12_io_in_valid_0),
    .io_in_valid_1(mesh_12_12_io_in_valid_1),
    .io_out_valid_0(mesh_12_12_io_out_valid_0),
    .io_out_valid_1(mesh_12_12_io_out_valid_1)
  );
  Tile mesh_12_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_13_clock),
    .io_in_a_0(mesh_12_13_io_in_a_0),
    .io_in_a_1(mesh_12_13_io_in_a_1),
    .io_in_b_0(mesh_12_13_io_in_b_0),
    .io_in_b_1(mesh_12_13_io_in_b_1),
    .io_in_d_0(mesh_12_13_io_in_d_0),
    .io_in_d_1(mesh_12_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_13_io_in_control_1_shift),
    .io_in_id_0(mesh_12_13_io_in_id_0),
    .io_in_id_1(mesh_12_13_io_in_id_1),
    .io_in_last_0(mesh_12_13_io_in_last_0),
    .io_in_last_1(mesh_12_13_io_in_last_1),
    .io_out_a_0(mesh_12_13_io_out_a_0),
    .io_out_a_1(mesh_12_13_io_out_a_1),
    .io_out_c_0(mesh_12_13_io_out_c_0),
    .io_out_c_1(mesh_12_13_io_out_c_1),
    .io_out_b_0(mesh_12_13_io_out_b_0),
    .io_out_b_1(mesh_12_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_13_io_out_control_1_shift),
    .io_out_id_0(mesh_12_13_io_out_id_0),
    .io_out_id_1(mesh_12_13_io_out_id_1),
    .io_out_last_0(mesh_12_13_io_out_last_0),
    .io_out_last_1(mesh_12_13_io_out_last_1),
    .io_in_valid_0(mesh_12_13_io_in_valid_0),
    .io_in_valid_1(mesh_12_13_io_in_valid_1),
    .io_out_valid_0(mesh_12_13_io_out_valid_0),
    .io_out_valid_1(mesh_12_13_io_out_valid_1)
  );
  Tile mesh_12_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_14_clock),
    .io_in_a_0(mesh_12_14_io_in_a_0),
    .io_in_a_1(mesh_12_14_io_in_a_1),
    .io_in_b_0(mesh_12_14_io_in_b_0),
    .io_in_b_1(mesh_12_14_io_in_b_1),
    .io_in_d_0(mesh_12_14_io_in_d_0),
    .io_in_d_1(mesh_12_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_14_io_in_control_1_shift),
    .io_in_id_0(mesh_12_14_io_in_id_0),
    .io_in_id_1(mesh_12_14_io_in_id_1),
    .io_in_last_0(mesh_12_14_io_in_last_0),
    .io_in_last_1(mesh_12_14_io_in_last_1),
    .io_out_a_0(mesh_12_14_io_out_a_0),
    .io_out_a_1(mesh_12_14_io_out_a_1),
    .io_out_c_0(mesh_12_14_io_out_c_0),
    .io_out_c_1(mesh_12_14_io_out_c_1),
    .io_out_b_0(mesh_12_14_io_out_b_0),
    .io_out_b_1(mesh_12_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_14_io_out_control_1_shift),
    .io_out_id_0(mesh_12_14_io_out_id_0),
    .io_out_id_1(mesh_12_14_io_out_id_1),
    .io_out_last_0(mesh_12_14_io_out_last_0),
    .io_out_last_1(mesh_12_14_io_out_last_1),
    .io_in_valid_0(mesh_12_14_io_in_valid_0),
    .io_in_valid_1(mesh_12_14_io_in_valid_1),
    .io_out_valid_0(mesh_12_14_io_out_valid_0),
    .io_out_valid_1(mesh_12_14_io_out_valid_1)
  );
  Tile mesh_12_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_12_15_clock),
    .io_in_a_0(mesh_12_15_io_in_a_0),
    .io_in_a_1(mesh_12_15_io_in_a_1),
    .io_in_b_0(mesh_12_15_io_in_b_0),
    .io_in_b_1(mesh_12_15_io_in_b_1),
    .io_in_d_0(mesh_12_15_io_in_d_0),
    .io_in_d_1(mesh_12_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_12_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_12_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_12_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_12_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_12_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_12_15_io_in_control_1_shift),
    .io_in_id_0(mesh_12_15_io_in_id_0),
    .io_in_id_1(mesh_12_15_io_in_id_1),
    .io_in_last_0(mesh_12_15_io_in_last_0),
    .io_in_last_1(mesh_12_15_io_in_last_1),
    .io_out_a_0(mesh_12_15_io_out_a_0),
    .io_out_a_1(mesh_12_15_io_out_a_1),
    .io_out_c_0(mesh_12_15_io_out_c_0),
    .io_out_c_1(mesh_12_15_io_out_c_1),
    .io_out_b_0(mesh_12_15_io_out_b_0),
    .io_out_b_1(mesh_12_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_12_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_12_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_12_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_12_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_12_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_12_15_io_out_control_1_shift),
    .io_out_id_0(mesh_12_15_io_out_id_0),
    .io_out_id_1(mesh_12_15_io_out_id_1),
    .io_out_last_0(mesh_12_15_io_out_last_0),
    .io_out_last_1(mesh_12_15_io_out_last_1),
    .io_in_valid_0(mesh_12_15_io_in_valid_0),
    .io_in_valid_1(mesh_12_15_io_in_valid_1),
    .io_out_valid_0(mesh_12_15_io_out_valid_0),
    .io_out_valid_1(mesh_12_15_io_out_valid_1)
  );
  Tile mesh_13_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_0_clock),
    .io_in_a_0(mesh_13_0_io_in_a_0),
    .io_in_a_1(mesh_13_0_io_in_a_1),
    .io_in_b_0(mesh_13_0_io_in_b_0),
    .io_in_b_1(mesh_13_0_io_in_b_1),
    .io_in_d_0(mesh_13_0_io_in_d_0),
    .io_in_d_1(mesh_13_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_0_io_in_control_1_shift),
    .io_in_id_0(mesh_13_0_io_in_id_0),
    .io_in_id_1(mesh_13_0_io_in_id_1),
    .io_in_last_0(mesh_13_0_io_in_last_0),
    .io_in_last_1(mesh_13_0_io_in_last_1),
    .io_out_a_0(mesh_13_0_io_out_a_0),
    .io_out_a_1(mesh_13_0_io_out_a_1),
    .io_out_c_0(mesh_13_0_io_out_c_0),
    .io_out_c_1(mesh_13_0_io_out_c_1),
    .io_out_b_0(mesh_13_0_io_out_b_0),
    .io_out_b_1(mesh_13_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_0_io_out_control_1_shift),
    .io_out_id_0(mesh_13_0_io_out_id_0),
    .io_out_id_1(mesh_13_0_io_out_id_1),
    .io_out_last_0(mesh_13_0_io_out_last_0),
    .io_out_last_1(mesh_13_0_io_out_last_1),
    .io_in_valid_0(mesh_13_0_io_in_valid_0),
    .io_in_valid_1(mesh_13_0_io_in_valid_1),
    .io_out_valid_0(mesh_13_0_io_out_valid_0),
    .io_out_valid_1(mesh_13_0_io_out_valid_1)
  );
  Tile mesh_13_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_1_clock),
    .io_in_a_0(mesh_13_1_io_in_a_0),
    .io_in_a_1(mesh_13_1_io_in_a_1),
    .io_in_b_0(mesh_13_1_io_in_b_0),
    .io_in_b_1(mesh_13_1_io_in_b_1),
    .io_in_d_0(mesh_13_1_io_in_d_0),
    .io_in_d_1(mesh_13_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_1_io_in_control_1_shift),
    .io_in_id_0(mesh_13_1_io_in_id_0),
    .io_in_id_1(mesh_13_1_io_in_id_1),
    .io_in_last_0(mesh_13_1_io_in_last_0),
    .io_in_last_1(mesh_13_1_io_in_last_1),
    .io_out_a_0(mesh_13_1_io_out_a_0),
    .io_out_a_1(mesh_13_1_io_out_a_1),
    .io_out_c_0(mesh_13_1_io_out_c_0),
    .io_out_c_1(mesh_13_1_io_out_c_1),
    .io_out_b_0(mesh_13_1_io_out_b_0),
    .io_out_b_1(mesh_13_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_1_io_out_control_1_shift),
    .io_out_id_0(mesh_13_1_io_out_id_0),
    .io_out_id_1(mesh_13_1_io_out_id_1),
    .io_out_last_0(mesh_13_1_io_out_last_0),
    .io_out_last_1(mesh_13_1_io_out_last_1),
    .io_in_valid_0(mesh_13_1_io_in_valid_0),
    .io_in_valid_1(mesh_13_1_io_in_valid_1),
    .io_out_valid_0(mesh_13_1_io_out_valid_0),
    .io_out_valid_1(mesh_13_1_io_out_valid_1)
  );
  Tile mesh_13_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_2_clock),
    .io_in_a_0(mesh_13_2_io_in_a_0),
    .io_in_a_1(mesh_13_2_io_in_a_1),
    .io_in_b_0(mesh_13_2_io_in_b_0),
    .io_in_b_1(mesh_13_2_io_in_b_1),
    .io_in_d_0(mesh_13_2_io_in_d_0),
    .io_in_d_1(mesh_13_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_2_io_in_control_1_shift),
    .io_in_id_0(mesh_13_2_io_in_id_0),
    .io_in_id_1(mesh_13_2_io_in_id_1),
    .io_in_last_0(mesh_13_2_io_in_last_0),
    .io_in_last_1(mesh_13_2_io_in_last_1),
    .io_out_a_0(mesh_13_2_io_out_a_0),
    .io_out_a_1(mesh_13_2_io_out_a_1),
    .io_out_c_0(mesh_13_2_io_out_c_0),
    .io_out_c_1(mesh_13_2_io_out_c_1),
    .io_out_b_0(mesh_13_2_io_out_b_0),
    .io_out_b_1(mesh_13_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_2_io_out_control_1_shift),
    .io_out_id_0(mesh_13_2_io_out_id_0),
    .io_out_id_1(mesh_13_2_io_out_id_1),
    .io_out_last_0(mesh_13_2_io_out_last_0),
    .io_out_last_1(mesh_13_2_io_out_last_1),
    .io_in_valid_0(mesh_13_2_io_in_valid_0),
    .io_in_valid_1(mesh_13_2_io_in_valid_1),
    .io_out_valid_0(mesh_13_2_io_out_valid_0),
    .io_out_valid_1(mesh_13_2_io_out_valid_1)
  );
  Tile mesh_13_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_3_clock),
    .io_in_a_0(mesh_13_3_io_in_a_0),
    .io_in_a_1(mesh_13_3_io_in_a_1),
    .io_in_b_0(mesh_13_3_io_in_b_0),
    .io_in_b_1(mesh_13_3_io_in_b_1),
    .io_in_d_0(mesh_13_3_io_in_d_0),
    .io_in_d_1(mesh_13_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_3_io_in_control_1_shift),
    .io_in_id_0(mesh_13_3_io_in_id_0),
    .io_in_id_1(mesh_13_3_io_in_id_1),
    .io_in_last_0(mesh_13_3_io_in_last_0),
    .io_in_last_1(mesh_13_3_io_in_last_1),
    .io_out_a_0(mesh_13_3_io_out_a_0),
    .io_out_a_1(mesh_13_3_io_out_a_1),
    .io_out_c_0(mesh_13_3_io_out_c_0),
    .io_out_c_1(mesh_13_3_io_out_c_1),
    .io_out_b_0(mesh_13_3_io_out_b_0),
    .io_out_b_1(mesh_13_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_3_io_out_control_1_shift),
    .io_out_id_0(mesh_13_3_io_out_id_0),
    .io_out_id_1(mesh_13_3_io_out_id_1),
    .io_out_last_0(mesh_13_3_io_out_last_0),
    .io_out_last_1(mesh_13_3_io_out_last_1),
    .io_in_valid_0(mesh_13_3_io_in_valid_0),
    .io_in_valid_1(mesh_13_3_io_in_valid_1),
    .io_out_valid_0(mesh_13_3_io_out_valid_0),
    .io_out_valid_1(mesh_13_3_io_out_valid_1)
  );
  Tile mesh_13_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_4_clock),
    .io_in_a_0(mesh_13_4_io_in_a_0),
    .io_in_a_1(mesh_13_4_io_in_a_1),
    .io_in_b_0(mesh_13_4_io_in_b_0),
    .io_in_b_1(mesh_13_4_io_in_b_1),
    .io_in_d_0(mesh_13_4_io_in_d_0),
    .io_in_d_1(mesh_13_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_4_io_in_control_1_shift),
    .io_in_id_0(mesh_13_4_io_in_id_0),
    .io_in_id_1(mesh_13_4_io_in_id_1),
    .io_in_last_0(mesh_13_4_io_in_last_0),
    .io_in_last_1(mesh_13_4_io_in_last_1),
    .io_out_a_0(mesh_13_4_io_out_a_0),
    .io_out_a_1(mesh_13_4_io_out_a_1),
    .io_out_c_0(mesh_13_4_io_out_c_0),
    .io_out_c_1(mesh_13_4_io_out_c_1),
    .io_out_b_0(mesh_13_4_io_out_b_0),
    .io_out_b_1(mesh_13_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_4_io_out_control_1_shift),
    .io_out_id_0(mesh_13_4_io_out_id_0),
    .io_out_id_1(mesh_13_4_io_out_id_1),
    .io_out_last_0(mesh_13_4_io_out_last_0),
    .io_out_last_1(mesh_13_4_io_out_last_1),
    .io_in_valid_0(mesh_13_4_io_in_valid_0),
    .io_in_valid_1(mesh_13_4_io_in_valid_1),
    .io_out_valid_0(mesh_13_4_io_out_valid_0),
    .io_out_valid_1(mesh_13_4_io_out_valid_1)
  );
  Tile mesh_13_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_5_clock),
    .io_in_a_0(mesh_13_5_io_in_a_0),
    .io_in_a_1(mesh_13_5_io_in_a_1),
    .io_in_b_0(mesh_13_5_io_in_b_0),
    .io_in_b_1(mesh_13_5_io_in_b_1),
    .io_in_d_0(mesh_13_5_io_in_d_0),
    .io_in_d_1(mesh_13_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_5_io_in_control_1_shift),
    .io_in_id_0(mesh_13_5_io_in_id_0),
    .io_in_id_1(mesh_13_5_io_in_id_1),
    .io_in_last_0(mesh_13_5_io_in_last_0),
    .io_in_last_1(mesh_13_5_io_in_last_1),
    .io_out_a_0(mesh_13_5_io_out_a_0),
    .io_out_a_1(mesh_13_5_io_out_a_1),
    .io_out_c_0(mesh_13_5_io_out_c_0),
    .io_out_c_1(mesh_13_5_io_out_c_1),
    .io_out_b_0(mesh_13_5_io_out_b_0),
    .io_out_b_1(mesh_13_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_5_io_out_control_1_shift),
    .io_out_id_0(mesh_13_5_io_out_id_0),
    .io_out_id_1(mesh_13_5_io_out_id_1),
    .io_out_last_0(mesh_13_5_io_out_last_0),
    .io_out_last_1(mesh_13_5_io_out_last_1),
    .io_in_valid_0(mesh_13_5_io_in_valid_0),
    .io_in_valid_1(mesh_13_5_io_in_valid_1),
    .io_out_valid_0(mesh_13_5_io_out_valid_0),
    .io_out_valid_1(mesh_13_5_io_out_valid_1)
  );
  Tile mesh_13_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_6_clock),
    .io_in_a_0(mesh_13_6_io_in_a_0),
    .io_in_a_1(mesh_13_6_io_in_a_1),
    .io_in_b_0(mesh_13_6_io_in_b_0),
    .io_in_b_1(mesh_13_6_io_in_b_1),
    .io_in_d_0(mesh_13_6_io_in_d_0),
    .io_in_d_1(mesh_13_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_6_io_in_control_1_shift),
    .io_in_id_0(mesh_13_6_io_in_id_0),
    .io_in_id_1(mesh_13_6_io_in_id_1),
    .io_in_last_0(mesh_13_6_io_in_last_0),
    .io_in_last_1(mesh_13_6_io_in_last_1),
    .io_out_a_0(mesh_13_6_io_out_a_0),
    .io_out_a_1(mesh_13_6_io_out_a_1),
    .io_out_c_0(mesh_13_6_io_out_c_0),
    .io_out_c_1(mesh_13_6_io_out_c_1),
    .io_out_b_0(mesh_13_6_io_out_b_0),
    .io_out_b_1(mesh_13_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_6_io_out_control_1_shift),
    .io_out_id_0(mesh_13_6_io_out_id_0),
    .io_out_id_1(mesh_13_6_io_out_id_1),
    .io_out_last_0(mesh_13_6_io_out_last_0),
    .io_out_last_1(mesh_13_6_io_out_last_1),
    .io_in_valid_0(mesh_13_6_io_in_valid_0),
    .io_in_valid_1(mesh_13_6_io_in_valid_1),
    .io_out_valid_0(mesh_13_6_io_out_valid_0),
    .io_out_valid_1(mesh_13_6_io_out_valid_1)
  );
  Tile mesh_13_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_7_clock),
    .io_in_a_0(mesh_13_7_io_in_a_0),
    .io_in_a_1(mesh_13_7_io_in_a_1),
    .io_in_b_0(mesh_13_7_io_in_b_0),
    .io_in_b_1(mesh_13_7_io_in_b_1),
    .io_in_d_0(mesh_13_7_io_in_d_0),
    .io_in_d_1(mesh_13_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_7_io_in_control_1_shift),
    .io_in_id_0(mesh_13_7_io_in_id_0),
    .io_in_id_1(mesh_13_7_io_in_id_1),
    .io_in_last_0(mesh_13_7_io_in_last_0),
    .io_in_last_1(mesh_13_7_io_in_last_1),
    .io_out_a_0(mesh_13_7_io_out_a_0),
    .io_out_a_1(mesh_13_7_io_out_a_1),
    .io_out_c_0(mesh_13_7_io_out_c_0),
    .io_out_c_1(mesh_13_7_io_out_c_1),
    .io_out_b_0(mesh_13_7_io_out_b_0),
    .io_out_b_1(mesh_13_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_7_io_out_control_1_shift),
    .io_out_id_0(mesh_13_7_io_out_id_0),
    .io_out_id_1(mesh_13_7_io_out_id_1),
    .io_out_last_0(mesh_13_7_io_out_last_0),
    .io_out_last_1(mesh_13_7_io_out_last_1),
    .io_in_valid_0(mesh_13_7_io_in_valid_0),
    .io_in_valid_1(mesh_13_7_io_in_valid_1),
    .io_out_valid_0(mesh_13_7_io_out_valid_0),
    .io_out_valid_1(mesh_13_7_io_out_valid_1)
  );
  Tile mesh_13_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_8_clock),
    .io_in_a_0(mesh_13_8_io_in_a_0),
    .io_in_a_1(mesh_13_8_io_in_a_1),
    .io_in_b_0(mesh_13_8_io_in_b_0),
    .io_in_b_1(mesh_13_8_io_in_b_1),
    .io_in_d_0(mesh_13_8_io_in_d_0),
    .io_in_d_1(mesh_13_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_8_io_in_control_1_shift),
    .io_in_id_0(mesh_13_8_io_in_id_0),
    .io_in_id_1(mesh_13_8_io_in_id_1),
    .io_in_last_0(mesh_13_8_io_in_last_0),
    .io_in_last_1(mesh_13_8_io_in_last_1),
    .io_out_a_0(mesh_13_8_io_out_a_0),
    .io_out_a_1(mesh_13_8_io_out_a_1),
    .io_out_c_0(mesh_13_8_io_out_c_0),
    .io_out_c_1(mesh_13_8_io_out_c_1),
    .io_out_b_0(mesh_13_8_io_out_b_0),
    .io_out_b_1(mesh_13_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_8_io_out_control_1_shift),
    .io_out_id_0(mesh_13_8_io_out_id_0),
    .io_out_id_1(mesh_13_8_io_out_id_1),
    .io_out_last_0(mesh_13_8_io_out_last_0),
    .io_out_last_1(mesh_13_8_io_out_last_1),
    .io_in_valid_0(mesh_13_8_io_in_valid_0),
    .io_in_valid_1(mesh_13_8_io_in_valid_1),
    .io_out_valid_0(mesh_13_8_io_out_valid_0),
    .io_out_valid_1(mesh_13_8_io_out_valid_1)
  );
  Tile mesh_13_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_9_clock),
    .io_in_a_0(mesh_13_9_io_in_a_0),
    .io_in_a_1(mesh_13_9_io_in_a_1),
    .io_in_b_0(mesh_13_9_io_in_b_0),
    .io_in_b_1(mesh_13_9_io_in_b_1),
    .io_in_d_0(mesh_13_9_io_in_d_0),
    .io_in_d_1(mesh_13_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_9_io_in_control_1_shift),
    .io_in_id_0(mesh_13_9_io_in_id_0),
    .io_in_id_1(mesh_13_9_io_in_id_1),
    .io_in_last_0(mesh_13_9_io_in_last_0),
    .io_in_last_1(mesh_13_9_io_in_last_1),
    .io_out_a_0(mesh_13_9_io_out_a_0),
    .io_out_a_1(mesh_13_9_io_out_a_1),
    .io_out_c_0(mesh_13_9_io_out_c_0),
    .io_out_c_1(mesh_13_9_io_out_c_1),
    .io_out_b_0(mesh_13_9_io_out_b_0),
    .io_out_b_1(mesh_13_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_9_io_out_control_1_shift),
    .io_out_id_0(mesh_13_9_io_out_id_0),
    .io_out_id_1(mesh_13_9_io_out_id_1),
    .io_out_last_0(mesh_13_9_io_out_last_0),
    .io_out_last_1(mesh_13_9_io_out_last_1),
    .io_in_valid_0(mesh_13_9_io_in_valid_0),
    .io_in_valid_1(mesh_13_9_io_in_valid_1),
    .io_out_valid_0(mesh_13_9_io_out_valid_0),
    .io_out_valid_1(mesh_13_9_io_out_valid_1)
  );
  Tile mesh_13_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_10_clock),
    .io_in_a_0(mesh_13_10_io_in_a_0),
    .io_in_a_1(mesh_13_10_io_in_a_1),
    .io_in_b_0(mesh_13_10_io_in_b_0),
    .io_in_b_1(mesh_13_10_io_in_b_1),
    .io_in_d_0(mesh_13_10_io_in_d_0),
    .io_in_d_1(mesh_13_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_10_io_in_control_1_shift),
    .io_in_id_0(mesh_13_10_io_in_id_0),
    .io_in_id_1(mesh_13_10_io_in_id_1),
    .io_in_last_0(mesh_13_10_io_in_last_0),
    .io_in_last_1(mesh_13_10_io_in_last_1),
    .io_out_a_0(mesh_13_10_io_out_a_0),
    .io_out_a_1(mesh_13_10_io_out_a_1),
    .io_out_c_0(mesh_13_10_io_out_c_0),
    .io_out_c_1(mesh_13_10_io_out_c_1),
    .io_out_b_0(mesh_13_10_io_out_b_0),
    .io_out_b_1(mesh_13_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_10_io_out_control_1_shift),
    .io_out_id_0(mesh_13_10_io_out_id_0),
    .io_out_id_1(mesh_13_10_io_out_id_1),
    .io_out_last_0(mesh_13_10_io_out_last_0),
    .io_out_last_1(mesh_13_10_io_out_last_1),
    .io_in_valid_0(mesh_13_10_io_in_valid_0),
    .io_in_valid_1(mesh_13_10_io_in_valid_1),
    .io_out_valid_0(mesh_13_10_io_out_valid_0),
    .io_out_valid_1(mesh_13_10_io_out_valid_1)
  );
  Tile mesh_13_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_11_clock),
    .io_in_a_0(mesh_13_11_io_in_a_0),
    .io_in_a_1(mesh_13_11_io_in_a_1),
    .io_in_b_0(mesh_13_11_io_in_b_0),
    .io_in_b_1(mesh_13_11_io_in_b_1),
    .io_in_d_0(mesh_13_11_io_in_d_0),
    .io_in_d_1(mesh_13_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_11_io_in_control_1_shift),
    .io_in_id_0(mesh_13_11_io_in_id_0),
    .io_in_id_1(mesh_13_11_io_in_id_1),
    .io_in_last_0(mesh_13_11_io_in_last_0),
    .io_in_last_1(mesh_13_11_io_in_last_1),
    .io_out_a_0(mesh_13_11_io_out_a_0),
    .io_out_a_1(mesh_13_11_io_out_a_1),
    .io_out_c_0(mesh_13_11_io_out_c_0),
    .io_out_c_1(mesh_13_11_io_out_c_1),
    .io_out_b_0(mesh_13_11_io_out_b_0),
    .io_out_b_1(mesh_13_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_11_io_out_control_1_shift),
    .io_out_id_0(mesh_13_11_io_out_id_0),
    .io_out_id_1(mesh_13_11_io_out_id_1),
    .io_out_last_0(mesh_13_11_io_out_last_0),
    .io_out_last_1(mesh_13_11_io_out_last_1),
    .io_in_valid_0(mesh_13_11_io_in_valid_0),
    .io_in_valid_1(mesh_13_11_io_in_valid_1),
    .io_out_valid_0(mesh_13_11_io_out_valid_0),
    .io_out_valid_1(mesh_13_11_io_out_valid_1)
  );
  Tile mesh_13_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_12_clock),
    .io_in_a_0(mesh_13_12_io_in_a_0),
    .io_in_a_1(mesh_13_12_io_in_a_1),
    .io_in_b_0(mesh_13_12_io_in_b_0),
    .io_in_b_1(mesh_13_12_io_in_b_1),
    .io_in_d_0(mesh_13_12_io_in_d_0),
    .io_in_d_1(mesh_13_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_12_io_in_control_1_shift),
    .io_in_id_0(mesh_13_12_io_in_id_0),
    .io_in_id_1(mesh_13_12_io_in_id_1),
    .io_in_last_0(mesh_13_12_io_in_last_0),
    .io_in_last_1(mesh_13_12_io_in_last_1),
    .io_out_a_0(mesh_13_12_io_out_a_0),
    .io_out_a_1(mesh_13_12_io_out_a_1),
    .io_out_c_0(mesh_13_12_io_out_c_0),
    .io_out_c_1(mesh_13_12_io_out_c_1),
    .io_out_b_0(mesh_13_12_io_out_b_0),
    .io_out_b_1(mesh_13_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_12_io_out_control_1_shift),
    .io_out_id_0(mesh_13_12_io_out_id_0),
    .io_out_id_1(mesh_13_12_io_out_id_1),
    .io_out_last_0(mesh_13_12_io_out_last_0),
    .io_out_last_1(mesh_13_12_io_out_last_1),
    .io_in_valid_0(mesh_13_12_io_in_valid_0),
    .io_in_valid_1(mesh_13_12_io_in_valid_1),
    .io_out_valid_0(mesh_13_12_io_out_valid_0),
    .io_out_valid_1(mesh_13_12_io_out_valid_1)
  );
  Tile mesh_13_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_13_clock),
    .io_in_a_0(mesh_13_13_io_in_a_0),
    .io_in_a_1(mesh_13_13_io_in_a_1),
    .io_in_b_0(mesh_13_13_io_in_b_0),
    .io_in_b_1(mesh_13_13_io_in_b_1),
    .io_in_d_0(mesh_13_13_io_in_d_0),
    .io_in_d_1(mesh_13_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_13_io_in_control_1_shift),
    .io_in_id_0(mesh_13_13_io_in_id_0),
    .io_in_id_1(mesh_13_13_io_in_id_1),
    .io_in_last_0(mesh_13_13_io_in_last_0),
    .io_in_last_1(mesh_13_13_io_in_last_1),
    .io_out_a_0(mesh_13_13_io_out_a_0),
    .io_out_a_1(mesh_13_13_io_out_a_1),
    .io_out_c_0(mesh_13_13_io_out_c_0),
    .io_out_c_1(mesh_13_13_io_out_c_1),
    .io_out_b_0(mesh_13_13_io_out_b_0),
    .io_out_b_1(mesh_13_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_13_io_out_control_1_shift),
    .io_out_id_0(mesh_13_13_io_out_id_0),
    .io_out_id_1(mesh_13_13_io_out_id_1),
    .io_out_last_0(mesh_13_13_io_out_last_0),
    .io_out_last_1(mesh_13_13_io_out_last_1),
    .io_in_valid_0(mesh_13_13_io_in_valid_0),
    .io_in_valid_1(mesh_13_13_io_in_valid_1),
    .io_out_valid_0(mesh_13_13_io_out_valid_0),
    .io_out_valid_1(mesh_13_13_io_out_valid_1)
  );
  Tile mesh_13_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_14_clock),
    .io_in_a_0(mesh_13_14_io_in_a_0),
    .io_in_a_1(mesh_13_14_io_in_a_1),
    .io_in_b_0(mesh_13_14_io_in_b_0),
    .io_in_b_1(mesh_13_14_io_in_b_1),
    .io_in_d_0(mesh_13_14_io_in_d_0),
    .io_in_d_1(mesh_13_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_14_io_in_control_1_shift),
    .io_in_id_0(mesh_13_14_io_in_id_0),
    .io_in_id_1(mesh_13_14_io_in_id_1),
    .io_in_last_0(mesh_13_14_io_in_last_0),
    .io_in_last_1(mesh_13_14_io_in_last_1),
    .io_out_a_0(mesh_13_14_io_out_a_0),
    .io_out_a_1(mesh_13_14_io_out_a_1),
    .io_out_c_0(mesh_13_14_io_out_c_0),
    .io_out_c_1(mesh_13_14_io_out_c_1),
    .io_out_b_0(mesh_13_14_io_out_b_0),
    .io_out_b_1(mesh_13_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_14_io_out_control_1_shift),
    .io_out_id_0(mesh_13_14_io_out_id_0),
    .io_out_id_1(mesh_13_14_io_out_id_1),
    .io_out_last_0(mesh_13_14_io_out_last_0),
    .io_out_last_1(mesh_13_14_io_out_last_1),
    .io_in_valid_0(mesh_13_14_io_in_valid_0),
    .io_in_valid_1(mesh_13_14_io_in_valid_1),
    .io_out_valid_0(mesh_13_14_io_out_valid_0),
    .io_out_valid_1(mesh_13_14_io_out_valid_1)
  );
  Tile mesh_13_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_13_15_clock),
    .io_in_a_0(mesh_13_15_io_in_a_0),
    .io_in_a_1(mesh_13_15_io_in_a_1),
    .io_in_b_0(mesh_13_15_io_in_b_0),
    .io_in_b_1(mesh_13_15_io_in_b_1),
    .io_in_d_0(mesh_13_15_io_in_d_0),
    .io_in_d_1(mesh_13_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_13_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_13_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_13_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_13_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_13_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_13_15_io_in_control_1_shift),
    .io_in_id_0(mesh_13_15_io_in_id_0),
    .io_in_id_1(mesh_13_15_io_in_id_1),
    .io_in_last_0(mesh_13_15_io_in_last_0),
    .io_in_last_1(mesh_13_15_io_in_last_1),
    .io_out_a_0(mesh_13_15_io_out_a_0),
    .io_out_a_1(mesh_13_15_io_out_a_1),
    .io_out_c_0(mesh_13_15_io_out_c_0),
    .io_out_c_1(mesh_13_15_io_out_c_1),
    .io_out_b_0(mesh_13_15_io_out_b_0),
    .io_out_b_1(mesh_13_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_13_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_13_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_13_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_13_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_13_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_13_15_io_out_control_1_shift),
    .io_out_id_0(mesh_13_15_io_out_id_0),
    .io_out_id_1(mesh_13_15_io_out_id_1),
    .io_out_last_0(mesh_13_15_io_out_last_0),
    .io_out_last_1(mesh_13_15_io_out_last_1),
    .io_in_valid_0(mesh_13_15_io_in_valid_0),
    .io_in_valid_1(mesh_13_15_io_in_valid_1),
    .io_out_valid_0(mesh_13_15_io_out_valid_0),
    .io_out_valid_1(mesh_13_15_io_out_valid_1)
  );
  Tile mesh_14_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_0_clock),
    .io_in_a_0(mesh_14_0_io_in_a_0),
    .io_in_a_1(mesh_14_0_io_in_a_1),
    .io_in_b_0(mesh_14_0_io_in_b_0),
    .io_in_b_1(mesh_14_0_io_in_b_1),
    .io_in_d_0(mesh_14_0_io_in_d_0),
    .io_in_d_1(mesh_14_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_0_io_in_control_1_shift),
    .io_in_id_0(mesh_14_0_io_in_id_0),
    .io_in_id_1(mesh_14_0_io_in_id_1),
    .io_in_last_0(mesh_14_0_io_in_last_0),
    .io_in_last_1(mesh_14_0_io_in_last_1),
    .io_out_a_0(mesh_14_0_io_out_a_0),
    .io_out_a_1(mesh_14_0_io_out_a_1),
    .io_out_c_0(mesh_14_0_io_out_c_0),
    .io_out_c_1(mesh_14_0_io_out_c_1),
    .io_out_b_0(mesh_14_0_io_out_b_0),
    .io_out_b_1(mesh_14_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_0_io_out_control_1_shift),
    .io_out_id_0(mesh_14_0_io_out_id_0),
    .io_out_id_1(mesh_14_0_io_out_id_1),
    .io_out_last_0(mesh_14_0_io_out_last_0),
    .io_out_last_1(mesh_14_0_io_out_last_1),
    .io_in_valid_0(mesh_14_0_io_in_valid_0),
    .io_in_valid_1(mesh_14_0_io_in_valid_1),
    .io_out_valid_0(mesh_14_0_io_out_valid_0),
    .io_out_valid_1(mesh_14_0_io_out_valid_1)
  );
  Tile mesh_14_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_1_clock),
    .io_in_a_0(mesh_14_1_io_in_a_0),
    .io_in_a_1(mesh_14_1_io_in_a_1),
    .io_in_b_0(mesh_14_1_io_in_b_0),
    .io_in_b_1(mesh_14_1_io_in_b_1),
    .io_in_d_0(mesh_14_1_io_in_d_0),
    .io_in_d_1(mesh_14_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_1_io_in_control_1_shift),
    .io_in_id_0(mesh_14_1_io_in_id_0),
    .io_in_id_1(mesh_14_1_io_in_id_1),
    .io_in_last_0(mesh_14_1_io_in_last_0),
    .io_in_last_1(mesh_14_1_io_in_last_1),
    .io_out_a_0(mesh_14_1_io_out_a_0),
    .io_out_a_1(mesh_14_1_io_out_a_1),
    .io_out_c_0(mesh_14_1_io_out_c_0),
    .io_out_c_1(mesh_14_1_io_out_c_1),
    .io_out_b_0(mesh_14_1_io_out_b_0),
    .io_out_b_1(mesh_14_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_1_io_out_control_1_shift),
    .io_out_id_0(mesh_14_1_io_out_id_0),
    .io_out_id_1(mesh_14_1_io_out_id_1),
    .io_out_last_0(mesh_14_1_io_out_last_0),
    .io_out_last_1(mesh_14_1_io_out_last_1),
    .io_in_valid_0(mesh_14_1_io_in_valid_0),
    .io_in_valid_1(mesh_14_1_io_in_valid_1),
    .io_out_valid_0(mesh_14_1_io_out_valid_0),
    .io_out_valid_1(mesh_14_1_io_out_valid_1)
  );
  Tile mesh_14_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_2_clock),
    .io_in_a_0(mesh_14_2_io_in_a_0),
    .io_in_a_1(mesh_14_2_io_in_a_1),
    .io_in_b_0(mesh_14_2_io_in_b_0),
    .io_in_b_1(mesh_14_2_io_in_b_1),
    .io_in_d_0(mesh_14_2_io_in_d_0),
    .io_in_d_1(mesh_14_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_2_io_in_control_1_shift),
    .io_in_id_0(mesh_14_2_io_in_id_0),
    .io_in_id_1(mesh_14_2_io_in_id_1),
    .io_in_last_0(mesh_14_2_io_in_last_0),
    .io_in_last_1(mesh_14_2_io_in_last_1),
    .io_out_a_0(mesh_14_2_io_out_a_0),
    .io_out_a_1(mesh_14_2_io_out_a_1),
    .io_out_c_0(mesh_14_2_io_out_c_0),
    .io_out_c_1(mesh_14_2_io_out_c_1),
    .io_out_b_0(mesh_14_2_io_out_b_0),
    .io_out_b_1(mesh_14_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_2_io_out_control_1_shift),
    .io_out_id_0(mesh_14_2_io_out_id_0),
    .io_out_id_1(mesh_14_2_io_out_id_1),
    .io_out_last_0(mesh_14_2_io_out_last_0),
    .io_out_last_1(mesh_14_2_io_out_last_1),
    .io_in_valid_0(mesh_14_2_io_in_valid_0),
    .io_in_valid_1(mesh_14_2_io_in_valid_1),
    .io_out_valid_0(mesh_14_2_io_out_valid_0),
    .io_out_valid_1(mesh_14_2_io_out_valid_1)
  );
  Tile mesh_14_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_3_clock),
    .io_in_a_0(mesh_14_3_io_in_a_0),
    .io_in_a_1(mesh_14_3_io_in_a_1),
    .io_in_b_0(mesh_14_3_io_in_b_0),
    .io_in_b_1(mesh_14_3_io_in_b_1),
    .io_in_d_0(mesh_14_3_io_in_d_0),
    .io_in_d_1(mesh_14_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_3_io_in_control_1_shift),
    .io_in_id_0(mesh_14_3_io_in_id_0),
    .io_in_id_1(mesh_14_3_io_in_id_1),
    .io_in_last_0(mesh_14_3_io_in_last_0),
    .io_in_last_1(mesh_14_3_io_in_last_1),
    .io_out_a_0(mesh_14_3_io_out_a_0),
    .io_out_a_1(mesh_14_3_io_out_a_1),
    .io_out_c_0(mesh_14_3_io_out_c_0),
    .io_out_c_1(mesh_14_3_io_out_c_1),
    .io_out_b_0(mesh_14_3_io_out_b_0),
    .io_out_b_1(mesh_14_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_3_io_out_control_1_shift),
    .io_out_id_0(mesh_14_3_io_out_id_0),
    .io_out_id_1(mesh_14_3_io_out_id_1),
    .io_out_last_0(mesh_14_3_io_out_last_0),
    .io_out_last_1(mesh_14_3_io_out_last_1),
    .io_in_valid_0(mesh_14_3_io_in_valid_0),
    .io_in_valid_1(mesh_14_3_io_in_valid_1),
    .io_out_valid_0(mesh_14_3_io_out_valid_0),
    .io_out_valid_1(mesh_14_3_io_out_valid_1)
  );
  Tile mesh_14_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_4_clock),
    .io_in_a_0(mesh_14_4_io_in_a_0),
    .io_in_a_1(mesh_14_4_io_in_a_1),
    .io_in_b_0(mesh_14_4_io_in_b_0),
    .io_in_b_1(mesh_14_4_io_in_b_1),
    .io_in_d_0(mesh_14_4_io_in_d_0),
    .io_in_d_1(mesh_14_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_4_io_in_control_1_shift),
    .io_in_id_0(mesh_14_4_io_in_id_0),
    .io_in_id_1(mesh_14_4_io_in_id_1),
    .io_in_last_0(mesh_14_4_io_in_last_0),
    .io_in_last_1(mesh_14_4_io_in_last_1),
    .io_out_a_0(mesh_14_4_io_out_a_0),
    .io_out_a_1(mesh_14_4_io_out_a_1),
    .io_out_c_0(mesh_14_4_io_out_c_0),
    .io_out_c_1(mesh_14_4_io_out_c_1),
    .io_out_b_0(mesh_14_4_io_out_b_0),
    .io_out_b_1(mesh_14_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_4_io_out_control_1_shift),
    .io_out_id_0(mesh_14_4_io_out_id_0),
    .io_out_id_1(mesh_14_4_io_out_id_1),
    .io_out_last_0(mesh_14_4_io_out_last_0),
    .io_out_last_1(mesh_14_4_io_out_last_1),
    .io_in_valid_0(mesh_14_4_io_in_valid_0),
    .io_in_valid_1(mesh_14_4_io_in_valid_1),
    .io_out_valid_0(mesh_14_4_io_out_valid_0),
    .io_out_valid_1(mesh_14_4_io_out_valid_1)
  );
  Tile mesh_14_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_5_clock),
    .io_in_a_0(mesh_14_5_io_in_a_0),
    .io_in_a_1(mesh_14_5_io_in_a_1),
    .io_in_b_0(mesh_14_5_io_in_b_0),
    .io_in_b_1(mesh_14_5_io_in_b_1),
    .io_in_d_0(mesh_14_5_io_in_d_0),
    .io_in_d_1(mesh_14_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_5_io_in_control_1_shift),
    .io_in_id_0(mesh_14_5_io_in_id_0),
    .io_in_id_1(mesh_14_5_io_in_id_1),
    .io_in_last_0(mesh_14_5_io_in_last_0),
    .io_in_last_1(mesh_14_5_io_in_last_1),
    .io_out_a_0(mesh_14_5_io_out_a_0),
    .io_out_a_1(mesh_14_5_io_out_a_1),
    .io_out_c_0(mesh_14_5_io_out_c_0),
    .io_out_c_1(mesh_14_5_io_out_c_1),
    .io_out_b_0(mesh_14_5_io_out_b_0),
    .io_out_b_1(mesh_14_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_5_io_out_control_1_shift),
    .io_out_id_0(mesh_14_5_io_out_id_0),
    .io_out_id_1(mesh_14_5_io_out_id_1),
    .io_out_last_0(mesh_14_5_io_out_last_0),
    .io_out_last_1(mesh_14_5_io_out_last_1),
    .io_in_valid_0(mesh_14_5_io_in_valid_0),
    .io_in_valid_1(mesh_14_5_io_in_valid_1),
    .io_out_valid_0(mesh_14_5_io_out_valid_0),
    .io_out_valid_1(mesh_14_5_io_out_valid_1)
  );
  Tile mesh_14_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_6_clock),
    .io_in_a_0(mesh_14_6_io_in_a_0),
    .io_in_a_1(mesh_14_6_io_in_a_1),
    .io_in_b_0(mesh_14_6_io_in_b_0),
    .io_in_b_1(mesh_14_6_io_in_b_1),
    .io_in_d_0(mesh_14_6_io_in_d_0),
    .io_in_d_1(mesh_14_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_6_io_in_control_1_shift),
    .io_in_id_0(mesh_14_6_io_in_id_0),
    .io_in_id_1(mesh_14_6_io_in_id_1),
    .io_in_last_0(mesh_14_6_io_in_last_0),
    .io_in_last_1(mesh_14_6_io_in_last_1),
    .io_out_a_0(mesh_14_6_io_out_a_0),
    .io_out_a_1(mesh_14_6_io_out_a_1),
    .io_out_c_0(mesh_14_6_io_out_c_0),
    .io_out_c_1(mesh_14_6_io_out_c_1),
    .io_out_b_0(mesh_14_6_io_out_b_0),
    .io_out_b_1(mesh_14_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_6_io_out_control_1_shift),
    .io_out_id_0(mesh_14_6_io_out_id_0),
    .io_out_id_1(mesh_14_6_io_out_id_1),
    .io_out_last_0(mesh_14_6_io_out_last_0),
    .io_out_last_1(mesh_14_6_io_out_last_1),
    .io_in_valid_0(mesh_14_6_io_in_valid_0),
    .io_in_valid_1(mesh_14_6_io_in_valid_1),
    .io_out_valid_0(mesh_14_6_io_out_valid_0),
    .io_out_valid_1(mesh_14_6_io_out_valid_1)
  );
  Tile mesh_14_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_7_clock),
    .io_in_a_0(mesh_14_7_io_in_a_0),
    .io_in_a_1(mesh_14_7_io_in_a_1),
    .io_in_b_0(mesh_14_7_io_in_b_0),
    .io_in_b_1(mesh_14_7_io_in_b_1),
    .io_in_d_0(mesh_14_7_io_in_d_0),
    .io_in_d_1(mesh_14_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_7_io_in_control_1_shift),
    .io_in_id_0(mesh_14_7_io_in_id_0),
    .io_in_id_1(mesh_14_7_io_in_id_1),
    .io_in_last_0(mesh_14_7_io_in_last_0),
    .io_in_last_1(mesh_14_7_io_in_last_1),
    .io_out_a_0(mesh_14_7_io_out_a_0),
    .io_out_a_1(mesh_14_7_io_out_a_1),
    .io_out_c_0(mesh_14_7_io_out_c_0),
    .io_out_c_1(mesh_14_7_io_out_c_1),
    .io_out_b_0(mesh_14_7_io_out_b_0),
    .io_out_b_1(mesh_14_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_7_io_out_control_1_shift),
    .io_out_id_0(mesh_14_7_io_out_id_0),
    .io_out_id_1(mesh_14_7_io_out_id_1),
    .io_out_last_0(mesh_14_7_io_out_last_0),
    .io_out_last_1(mesh_14_7_io_out_last_1),
    .io_in_valid_0(mesh_14_7_io_in_valid_0),
    .io_in_valid_1(mesh_14_7_io_in_valid_1),
    .io_out_valid_0(mesh_14_7_io_out_valid_0),
    .io_out_valid_1(mesh_14_7_io_out_valid_1)
  );
  Tile mesh_14_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_8_clock),
    .io_in_a_0(mesh_14_8_io_in_a_0),
    .io_in_a_1(mesh_14_8_io_in_a_1),
    .io_in_b_0(mesh_14_8_io_in_b_0),
    .io_in_b_1(mesh_14_8_io_in_b_1),
    .io_in_d_0(mesh_14_8_io_in_d_0),
    .io_in_d_1(mesh_14_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_8_io_in_control_1_shift),
    .io_in_id_0(mesh_14_8_io_in_id_0),
    .io_in_id_1(mesh_14_8_io_in_id_1),
    .io_in_last_0(mesh_14_8_io_in_last_0),
    .io_in_last_1(mesh_14_8_io_in_last_1),
    .io_out_a_0(mesh_14_8_io_out_a_0),
    .io_out_a_1(mesh_14_8_io_out_a_1),
    .io_out_c_0(mesh_14_8_io_out_c_0),
    .io_out_c_1(mesh_14_8_io_out_c_1),
    .io_out_b_0(mesh_14_8_io_out_b_0),
    .io_out_b_1(mesh_14_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_8_io_out_control_1_shift),
    .io_out_id_0(mesh_14_8_io_out_id_0),
    .io_out_id_1(mesh_14_8_io_out_id_1),
    .io_out_last_0(mesh_14_8_io_out_last_0),
    .io_out_last_1(mesh_14_8_io_out_last_1),
    .io_in_valid_0(mesh_14_8_io_in_valid_0),
    .io_in_valid_1(mesh_14_8_io_in_valid_1),
    .io_out_valid_0(mesh_14_8_io_out_valid_0),
    .io_out_valid_1(mesh_14_8_io_out_valid_1)
  );
  Tile mesh_14_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_9_clock),
    .io_in_a_0(mesh_14_9_io_in_a_0),
    .io_in_a_1(mesh_14_9_io_in_a_1),
    .io_in_b_0(mesh_14_9_io_in_b_0),
    .io_in_b_1(mesh_14_9_io_in_b_1),
    .io_in_d_0(mesh_14_9_io_in_d_0),
    .io_in_d_1(mesh_14_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_9_io_in_control_1_shift),
    .io_in_id_0(mesh_14_9_io_in_id_0),
    .io_in_id_1(mesh_14_9_io_in_id_1),
    .io_in_last_0(mesh_14_9_io_in_last_0),
    .io_in_last_1(mesh_14_9_io_in_last_1),
    .io_out_a_0(mesh_14_9_io_out_a_0),
    .io_out_a_1(mesh_14_9_io_out_a_1),
    .io_out_c_0(mesh_14_9_io_out_c_0),
    .io_out_c_1(mesh_14_9_io_out_c_1),
    .io_out_b_0(mesh_14_9_io_out_b_0),
    .io_out_b_1(mesh_14_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_9_io_out_control_1_shift),
    .io_out_id_0(mesh_14_9_io_out_id_0),
    .io_out_id_1(mesh_14_9_io_out_id_1),
    .io_out_last_0(mesh_14_9_io_out_last_0),
    .io_out_last_1(mesh_14_9_io_out_last_1),
    .io_in_valid_0(mesh_14_9_io_in_valid_0),
    .io_in_valid_1(mesh_14_9_io_in_valid_1),
    .io_out_valid_0(mesh_14_9_io_out_valid_0),
    .io_out_valid_1(mesh_14_9_io_out_valid_1)
  );
  Tile mesh_14_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_10_clock),
    .io_in_a_0(mesh_14_10_io_in_a_0),
    .io_in_a_1(mesh_14_10_io_in_a_1),
    .io_in_b_0(mesh_14_10_io_in_b_0),
    .io_in_b_1(mesh_14_10_io_in_b_1),
    .io_in_d_0(mesh_14_10_io_in_d_0),
    .io_in_d_1(mesh_14_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_10_io_in_control_1_shift),
    .io_in_id_0(mesh_14_10_io_in_id_0),
    .io_in_id_1(mesh_14_10_io_in_id_1),
    .io_in_last_0(mesh_14_10_io_in_last_0),
    .io_in_last_1(mesh_14_10_io_in_last_1),
    .io_out_a_0(mesh_14_10_io_out_a_0),
    .io_out_a_1(mesh_14_10_io_out_a_1),
    .io_out_c_0(mesh_14_10_io_out_c_0),
    .io_out_c_1(mesh_14_10_io_out_c_1),
    .io_out_b_0(mesh_14_10_io_out_b_0),
    .io_out_b_1(mesh_14_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_10_io_out_control_1_shift),
    .io_out_id_0(mesh_14_10_io_out_id_0),
    .io_out_id_1(mesh_14_10_io_out_id_1),
    .io_out_last_0(mesh_14_10_io_out_last_0),
    .io_out_last_1(mesh_14_10_io_out_last_1),
    .io_in_valid_0(mesh_14_10_io_in_valid_0),
    .io_in_valid_1(mesh_14_10_io_in_valid_1),
    .io_out_valid_0(mesh_14_10_io_out_valid_0),
    .io_out_valid_1(mesh_14_10_io_out_valid_1)
  );
  Tile mesh_14_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_11_clock),
    .io_in_a_0(mesh_14_11_io_in_a_0),
    .io_in_a_1(mesh_14_11_io_in_a_1),
    .io_in_b_0(mesh_14_11_io_in_b_0),
    .io_in_b_1(mesh_14_11_io_in_b_1),
    .io_in_d_0(mesh_14_11_io_in_d_0),
    .io_in_d_1(mesh_14_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_11_io_in_control_1_shift),
    .io_in_id_0(mesh_14_11_io_in_id_0),
    .io_in_id_1(mesh_14_11_io_in_id_1),
    .io_in_last_0(mesh_14_11_io_in_last_0),
    .io_in_last_1(mesh_14_11_io_in_last_1),
    .io_out_a_0(mesh_14_11_io_out_a_0),
    .io_out_a_1(mesh_14_11_io_out_a_1),
    .io_out_c_0(mesh_14_11_io_out_c_0),
    .io_out_c_1(mesh_14_11_io_out_c_1),
    .io_out_b_0(mesh_14_11_io_out_b_0),
    .io_out_b_1(mesh_14_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_11_io_out_control_1_shift),
    .io_out_id_0(mesh_14_11_io_out_id_0),
    .io_out_id_1(mesh_14_11_io_out_id_1),
    .io_out_last_0(mesh_14_11_io_out_last_0),
    .io_out_last_1(mesh_14_11_io_out_last_1),
    .io_in_valid_0(mesh_14_11_io_in_valid_0),
    .io_in_valid_1(mesh_14_11_io_in_valid_1),
    .io_out_valid_0(mesh_14_11_io_out_valid_0),
    .io_out_valid_1(mesh_14_11_io_out_valid_1)
  );
  Tile mesh_14_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_12_clock),
    .io_in_a_0(mesh_14_12_io_in_a_0),
    .io_in_a_1(mesh_14_12_io_in_a_1),
    .io_in_b_0(mesh_14_12_io_in_b_0),
    .io_in_b_1(mesh_14_12_io_in_b_1),
    .io_in_d_0(mesh_14_12_io_in_d_0),
    .io_in_d_1(mesh_14_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_12_io_in_control_1_shift),
    .io_in_id_0(mesh_14_12_io_in_id_0),
    .io_in_id_1(mesh_14_12_io_in_id_1),
    .io_in_last_0(mesh_14_12_io_in_last_0),
    .io_in_last_1(mesh_14_12_io_in_last_1),
    .io_out_a_0(mesh_14_12_io_out_a_0),
    .io_out_a_1(mesh_14_12_io_out_a_1),
    .io_out_c_0(mesh_14_12_io_out_c_0),
    .io_out_c_1(mesh_14_12_io_out_c_1),
    .io_out_b_0(mesh_14_12_io_out_b_0),
    .io_out_b_1(mesh_14_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_12_io_out_control_1_shift),
    .io_out_id_0(mesh_14_12_io_out_id_0),
    .io_out_id_1(mesh_14_12_io_out_id_1),
    .io_out_last_0(mesh_14_12_io_out_last_0),
    .io_out_last_1(mesh_14_12_io_out_last_1),
    .io_in_valid_0(mesh_14_12_io_in_valid_0),
    .io_in_valid_1(mesh_14_12_io_in_valid_1),
    .io_out_valid_0(mesh_14_12_io_out_valid_0),
    .io_out_valid_1(mesh_14_12_io_out_valid_1)
  );
  Tile mesh_14_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_13_clock),
    .io_in_a_0(mesh_14_13_io_in_a_0),
    .io_in_a_1(mesh_14_13_io_in_a_1),
    .io_in_b_0(mesh_14_13_io_in_b_0),
    .io_in_b_1(mesh_14_13_io_in_b_1),
    .io_in_d_0(mesh_14_13_io_in_d_0),
    .io_in_d_1(mesh_14_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_13_io_in_control_1_shift),
    .io_in_id_0(mesh_14_13_io_in_id_0),
    .io_in_id_1(mesh_14_13_io_in_id_1),
    .io_in_last_0(mesh_14_13_io_in_last_0),
    .io_in_last_1(mesh_14_13_io_in_last_1),
    .io_out_a_0(mesh_14_13_io_out_a_0),
    .io_out_a_1(mesh_14_13_io_out_a_1),
    .io_out_c_0(mesh_14_13_io_out_c_0),
    .io_out_c_1(mesh_14_13_io_out_c_1),
    .io_out_b_0(mesh_14_13_io_out_b_0),
    .io_out_b_1(mesh_14_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_13_io_out_control_1_shift),
    .io_out_id_0(mesh_14_13_io_out_id_0),
    .io_out_id_1(mesh_14_13_io_out_id_1),
    .io_out_last_0(mesh_14_13_io_out_last_0),
    .io_out_last_1(mesh_14_13_io_out_last_1),
    .io_in_valid_0(mesh_14_13_io_in_valid_0),
    .io_in_valid_1(mesh_14_13_io_in_valid_1),
    .io_out_valid_0(mesh_14_13_io_out_valid_0),
    .io_out_valid_1(mesh_14_13_io_out_valid_1)
  );
  Tile mesh_14_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_14_clock),
    .io_in_a_0(mesh_14_14_io_in_a_0),
    .io_in_a_1(mesh_14_14_io_in_a_1),
    .io_in_b_0(mesh_14_14_io_in_b_0),
    .io_in_b_1(mesh_14_14_io_in_b_1),
    .io_in_d_0(mesh_14_14_io_in_d_0),
    .io_in_d_1(mesh_14_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_14_io_in_control_1_shift),
    .io_in_id_0(mesh_14_14_io_in_id_0),
    .io_in_id_1(mesh_14_14_io_in_id_1),
    .io_in_last_0(mesh_14_14_io_in_last_0),
    .io_in_last_1(mesh_14_14_io_in_last_1),
    .io_out_a_0(mesh_14_14_io_out_a_0),
    .io_out_a_1(mesh_14_14_io_out_a_1),
    .io_out_c_0(mesh_14_14_io_out_c_0),
    .io_out_c_1(mesh_14_14_io_out_c_1),
    .io_out_b_0(mesh_14_14_io_out_b_0),
    .io_out_b_1(mesh_14_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_14_io_out_control_1_shift),
    .io_out_id_0(mesh_14_14_io_out_id_0),
    .io_out_id_1(mesh_14_14_io_out_id_1),
    .io_out_last_0(mesh_14_14_io_out_last_0),
    .io_out_last_1(mesh_14_14_io_out_last_1),
    .io_in_valid_0(mesh_14_14_io_in_valid_0),
    .io_in_valid_1(mesh_14_14_io_in_valid_1),
    .io_out_valid_0(mesh_14_14_io_out_valid_0),
    .io_out_valid_1(mesh_14_14_io_out_valid_1)
  );
  Tile mesh_14_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_14_15_clock),
    .io_in_a_0(mesh_14_15_io_in_a_0),
    .io_in_a_1(mesh_14_15_io_in_a_1),
    .io_in_b_0(mesh_14_15_io_in_b_0),
    .io_in_b_1(mesh_14_15_io_in_b_1),
    .io_in_d_0(mesh_14_15_io_in_d_0),
    .io_in_d_1(mesh_14_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_14_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_14_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_14_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_14_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_14_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_14_15_io_in_control_1_shift),
    .io_in_id_0(mesh_14_15_io_in_id_0),
    .io_in_id_1(mesh_14_15_io_in_id_1),
    .io_in_last_0(mesh_14_15_io_in_last_0),
    .io_in_last_1(mesh_14_15_io_in_last_1),
    .io_out_a_0(mesh_14_15_io_out_a_0),
    .io_out_a_1(mesh_14_15_io_out_a_1),
    .io_out_c_0(mesh_14_15_io_out_c_0),
    .io_out_c_1(mesh_14_15_io_out_c_1),
    .io_out_b_0(mesh_14_15_io_out_b_0),
    .io_out_b_1(mesh_14_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_14_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_14_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_14_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_14_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_14_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_14_15_io_out_control_1_shift),
    .io_out_id_0(mesh_14_15_io_out_id_0),
    .io_out_id_1(mesh_14_15_io_out_id_1),
    .io_out_last_0(mesh_14_15_io_out_last_0),
    .io_out_last_1(mesh_14_15_io_out_last_1),
    .io_in_valid_0(mesh_14_15_io_in_valid_0),
    .io_in_valid_1(mesh_14_15_io_in_valid_1),
    .io_out_valid_0(mesh_14_15_io_out_valid_0),
    .io_out_valid_1(mesh_14_15_io_out_valid_1)
  );
  Tile_240 mesh_15_0 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_0_clock),
    .io_in_a_0(mesh_15_0_io_in_a_0),
    .io_in_a_1(mesh_15_0_io_in_a_1),
    .io_in_b_0(mesh_15_0_io_in_b_0),
    .io_in_b_1(mesh_15_0_io_in_b_1),
    .io_in_d_0(mesh_15_0_io_in_d_0),
    .io_in_d_1(mesh_15_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_0_io_in_control_1_shift),
    .io_in_id_0(mesh_15_0_io_in_id_0),
    .io_in_id_1(mesh_15_0_io_in_id_1),
    .io_in_last_0(mesh_15_0_io_in_last_0),
    .io_in_last_1(mesh_15_0_io_in_last_1),
    .io_out_a_0(mesh_15_0_io_out_a_0),
    .io_out_a_1(mesh_15_0_io_out_a_1),
    .io_out_c_0(mesh_15_0_io_out_c_0),
    .io_out_c_1(mesh_15_0_io_out_c_1),
    .io_out_b_0(mesh_15_0_io_out_b_0),
    .io_out_b_1(mesh_15_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_0_io_out_control_1_shift),
    .io_out_id_0(mesh_15_0_io_out_id_0),
    .io_out_id_1(mesh_15_0_io_out_id_1),
    .io_out_last_0(mesh_15_0_io_out_last_0),
    .io_out_last_1(mesh_15_0_io_out_last_1),
    .io_in_valid_0(mesh_15_0_io_in_valid_0),
    .io_in_valid_1(mesh_15_0_io_in_valid_1),
    .io_out_valid_0(mesh_15_0_io_out_valid_0),
    .io_out_valid_1(mesh_15_0_io_out_valid_1)
  );
  Tile_240 mesh_15_1 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_1_clock),
    .io_in_a_0(mesh_15_1_io_in_a_0),
    .io_in_a_1(mesh_15_1_io_in_a_1),
    .io_in_b_0(mesh_15_1_io_in_b_0),
    .io_in_b_1(mesh_15_1_io_in_b_1),
    .io_in_d_0(mesh_15_1_io_in_d_0),
    .io_in_d_1(mesh_15_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_1_io_in_control_1_shift),
    .io_in_id_0(mesh_15_1_io_in_id_0),
    .io_in_id_1(mesh_15_1_io_in_id_1),
    .io_in_last_0(mesh_15_1_io_in_last_0),
    .io_in_last_1(mesh_15_1_io_in_last_1),
    .io_out_a_0(mesh_15_1_io_out_a_0),
    .io_out_a_1(mesh_15_1_io_out_a_1),
    .io_out_c_0(mesh_15_1_io_out_c_0),
    .io_out_c_1(mesh_15_1_io_out_c_1),
    .io_out_b_0(mesh_15_1_io_out_b_0),
    .io_out_b_1(mesh_15_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_1_io_out_control_1_shift),
    .io_out_id_0(mesh_15_1_io_out_id_0),
    .io_out_id_1(mesh_15_1_io_out_id_1),
    .io_out_last_0(mesh_15_1_io_out_last_0),
    .io_out_last_1(mesh_15_1_io_out_last_1),
    .io_in_valid_0(mesh_15_1_io_in_valid_0),
    .io_in_valid_1(mesh_15_1_io_in_valid_1),
    .io_out_valid_0(mesh_15_1_io_out_valid_0),
    .io_out_valid_1(mesh_15_1_io_out_valid_1)
  );
  Tile_240 mesh_15_2 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_2_clock),
    .io_in_a_0(mesh_15_2_io_in_a_0),
    .io_in_a_1(mesh_15_2_io_in_a_1),
    .io_in_b_0(mesh_15_2_io_in_b_0),
    .io_in_b_1(mesh_15_2_io_in_b_1),
    .io_in_d_0(mesh_15_2_io_in_d_0),
    .io_in_d_1(mesh_15_2_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_2_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_2_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_2_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_2_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_2_io_in_control_1_shift),
    .io_in_id_0(mesh_15_2_io_in_id_0),
    .io_in_id_1(mesh_15_2_io_in_id_1),
    .io_in_last_0(mesh_15_2_io_in_last_0),
    .io_in_last_1(mesh_15_2_io_in_last_1),
    .io_out_a_0(mesh_15_2_io_out_a_0),
    .io_out_a_1(mesh_15_2_io_out_a_1),
    .io_out_c_0(mesh_15_2_io_out_c_0),
    .io_out_c_1(mesh_15_2_io_out_c_1),
    .io_out_b_0(mesh_15_2_io_out_b_0),
    .io_out_b_1(mesh_15_2_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_2_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_2_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_2_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_2_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_2_io_out_control_1_shift),
    .io_out_id_0(mesh_15_2_io_out_id_0),
    .io_out_id_1(mesh_15_2_io_out_id_1),
    .io_out_last_0(mesh_15_2_io_out_last_0),
    .io_out_last_1(mesh_15_2_io_out_last_1),
    .io_in_valid_0(mesh_15_2_io_in_valid_0),
    .io_in_valid_1(mesh_15_2_io_in_valid_1),
    .io_out_valid_0(mesh_15_2_io_out_valid_0),
    .io_out_valid_1(mesh_15_2_io_out_valid_1)
  );
  Tile_240 mesh_15_3 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_3_clock),
    .io_in_a_0(mesh_15_3_io_in_a_0),
    .io_in_a_1(mesh_15_3_io_in_a_1),
    .io_in_b_0(mesh_15_3_io_in_b_0),
    .io_in_b_1(mesh_15_3_io_in_b_1),
    .io_in_d_0(mesh_15_3_io_in_d_0),
    .io_in_d_1(mesh_15_3_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_3_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_3_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_3_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_3_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_3_io_in_control_1_shift),
    .io_in_id_0(mesh_15_3_io_in_id_0),
    .io_in_id_1(mesh_15_3_io_in_id_1),
    .io_in_last_0(mesh_15_3_io_in_last_0),
    .io_in_last_1(mesh_15_3_io_in_last_1),
    .io_out_a_0(mesh_15_3_io_out_a_0),
    .io_out_a_1(mesh_15_3_io_out_a_1),
    .io_out_c_0(mesh_15_3_io_out_c_0),
    .io_out_c_1(mesh_15_3_io_out_c_1),
    .io_out_b_0(mesh_15_3_io_out_b_0),
    .io_out_b_1(mesh_15_3_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_3_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_3_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_3_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_3_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_3_io_out_control_1_shift),
    .io_out_id_0(mesh_15_3_io_out_id_0),
    .io_out_id_1(mesh_15_3_io_out_id_1),
    .io_out_last_0(mesh_15_3_io_out_last_0),
    .io_out_last_1(mesh_15_3_io_out_last_1),
    .io_in_valid_0(mesh_15_3_io_in_valid_0),
    .io_in_valid_1(mesh_15_3_io_in_valid_1),
    .io_out_valid_0(mesh_15_3_io_out_valid_0),
    .io_out_valid_1(mesh_15_3_io_out_valid_1)
  );
  Tile_240 mesh_15_4 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_4_clock),
    .io_in_a_0(mesh_15_4_io_in_a_0),
    .io_in_a_1(mesh_15_4_io_in_a_1),
    .io_in_b_0(mesh_15_4_io_in_b_0),
    .io_in_b_1(mesh_15_4_io_in_b_1),
    .io_in_d_0(mesh_15_4_io_in_d_0),
    .io_in_d_1(mesh_15_4_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_4_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_4_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_4_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_4_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_4_io_in_control_1_shift),
    .io_in_id_0(mesh_15_4_io_in_id_0),
    .io_in_id_1(mesh_15_4_io_in_id_1),
    .io_in_last_0(mesh_15_4_io_in_last_0),
    .io_in_last_1(mesh_15_4_io_in_last_1),
    .io_out_a_0(mesh_15_4_io_out_a_0),
    .io_out_a_1(mesh_15_4_io_out_a_1),
    .io_out_c_0(mesh_15_4_io_out_c_0),
    .io_out_c_1(mesh_15_4_io_out_c_1),
    .io_out_b_0(mesh_15_4_io_out_b_0),
    .io_out_b_1(mesh_15_4_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_4_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_4_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_4_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_4_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_4_io_out_control_1_shift),
    .io_out_id_0(mesh_15_4_io_out_id_0),
    .io_out_id_1(mesh_15_4_io_out_id_1),
    .io_out_last_0(mesh_15_4_io_out_last_0),
    .io_out_last_1(mesh_15_4_io_out_last_1),
    .io_in_valid_0(mesh_15_4_io_in_valid_0),
    .io_in_valid_1(mesh_15_4_io_in_valid_1),
    .io_out_valid_0(mesh_15_4_io_out_valid_0),
    .io_out_valid_1(mesh_15_4_io_out_valid_1)
  );
  Tile_240 mesh_15_5 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_5_clock),
    .io_in_a_0(mesh_15_5_io_in_a_0),
    .io_in_a_1(mesh_15_5_io_in_a_1),
    .io_in_b_0(mesh_15_5_io_in_b_0),
    .io_in_b_1(mesh_15_5_io_in_b_1),
    .io_in_d_0(mesh_15_5_io_in_d_0),
    .io_in_d_1(mesh_15_5_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_5_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_5_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_5_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_5_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_5_io_in_control_1_shift),
    .io_in_id_0(mesh_15_5_io_in_id_0),
    .io_in_id_1(mesh_15_5_io_in_id_1),
    .io_in_last_0(mesh_15_5_io_in_last_0),
    .io_in_last_1(mesh_15_5_io_in_last_1),
    .io_out_a_0(mesh_15_5_io_out_a_0),
    .io_out_a_1(mesh_15_5_io_out_a_1),
    .io_out_c_0(mesh_15_5_io_out_c_0),
    .io_out_c_1(mesh_15_5_io_out_c_1),
    .io_out_b_0(mesh_15_5_io_out_b_0),
    .io_out_b_1(mesh_15_5_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_5_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_5_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_5_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_5_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_5_io_out_control_1_shift),
    .io_out_id_0(mesh_15_5_io_out_id_0),
    .io_out_id_1(mesh_15_5_io_out_id_1),
    .io_out_last_0(mesh_15_5_io_out_last_0),
    .io_out_last_1(mesh_15_5_io_out_last_1),
    .io_in_valid_0(mesh_15_5_io_in_valid_0),
    .io_in_valid_1(mesh_15_5_io_in_valid_1),
    .io_out_valid_0(mesh_15_5_io_out_valid_0),
    .io_out_valid_1(mesh_15_5_io_out_valid_1)
  );
  Tile_240 mesh_15_6 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_6_clock),
    .io_in_a_0(mesh_15_6_io_in_a_0),
    .io_in_a_1(mesh_15_6_io_in_a_1),
    .io_in_b_0(mesh_15_6_io_in_b_0),
    .io_in_b_1(mesh_15_6_io_in_b_1),
    .io_in_d_0(mesh_15_6_io_in_d_0),
    .io_in_d_1(mesh_15_6_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_6_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_6_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_6_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_6_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_6_io_in_control_1_shift),
    .io_in_id_0(mesh_15_6_io_in_id_0),
    .io_in_id_1(mesh_15_6_io_in_id_1),
    .io_in_last_0(mesh_15_6_io_in_last_0),
    .io_in_last_1(mesh_15_6_io_in_last_1),
    .io_out_a_0(mesh_15_6_io_out_a_0),
    .io_out_a_1(mesh_15_6_io_out_a_1),
    .io_out_c_0(mesh_15_6_io_out_c_0),
    .io_out_c_1(mesh_15_6_io_out_c_1),
    .io_out_b_0(mesh_15_6_io_out_b_0),
    .io_out_b_1(mesh_15_6_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_6_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_6_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_6_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_6_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_6_io_out_control_1_shift),
    .io_out_id_0(mesh_15_6_io_out_id_0),
    .io_out_id_1(mesh_15_6_io_out_id_1),
    .io_out_last_0(mesh_15_6_io_out_last_0),
    .io_out_last_1(mesh_15_6_io_out_last_1),
    .io_in_valid_0(mesh_15_6_io_in_valid_0),
    .io_in_valid_1(mesh_15_6_io_in_valid_1),
    .io_out_valid_0(mesh_15_6_io_out_valid_0),
    .io_out_valid_1(mesh_15_6_io_out_valid_1)
  );
  Tile_240 mesh_15_7 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_7_clock),
    .io_in_a_0(mesh_15_7_io_in_a_0),
    .io_in_a_1(mesh_15_7_io_in_a_1),
    .io_in_b_0(mesh_15_7_io_in_b_0),
    .io_in_b_1(mesh_15_7_io_in_b_1),
    .io_in_d_0(mesh_15_7_io_in_d_0),
    .io_in_d_1(mesh_15_7_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_7_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_7_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_7_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_7_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_7_io_in_control_1_shift),
    .io_in_id_0(mesh_15_7_io_in_id_0),
    .io_in_id_1(mesh_15_7_io_in_id_1),
    .io_in_last_0(mesh_15_7_io_in_last_0),
    .io_in_last_1(mesh_15_7_io_in_last_1),
    .io_out_a_0(mesh_15_7_io_out_a_0),
    .io_out_a_1(mesh_15_7_io_out_a_1),
    .io_out_c_0(mesh_15_7_io_out_c_0),
    .io_out_c_1(mesh_15_7_io_out_c_1),
    .io_out_b_0(mesh_15_7_io_out_b_0),
    .io_out_b_1(mesh_15_7_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_7_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_7_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_7_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_7_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_7_io_out_control_1_shift),
    .io_out_id_0(mesh_15_7_io_out_id_0),
    .io_out_id_1(mesh_15_7_io_out_id_1),
    .io_out_last_0(mesh_15_7_io_out_last_0),
    .io_out_last_1(mesh_15_7_io_out_last_1),
    .io_in_valid_0(mesh_15_7_io_in_valid_0),
    .io_in_valid_1(mesh_15_7_io_in_valid_1),
    .io_out_valid_0(mesh_15_7_io_out_valid_0),
    .io_out_valid_1(mesh_15_7_io_out_valid_1)
  );
  Tile_240 mesh_15_8 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_8_clock),
    .io_in_a_0(mesh_15_8_io_in_a_0),
    .io_in_a_1(mesh_15_8_io_in_a_1),
    .io_in_b_0(mesh_15_8_io_in_b_0),
    .io_in_b_1(mesh_15_8_io_in_b_1),
    .io_in_d_0(mesh_15_8_io_in_d_0),
    .io_in_d_1(mesh_15_8_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_8_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_8_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_8_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_8_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_8_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_8_io_in_control_1_shift),
    .io_in_id_0(mesh_15_8_io_in_id_0),
    .io_in_id_1(mesh_15_8_io_in_id_1),
    .io_in_last_0(mesh_15_8_io_in_last_0),
    .io_in_last_1(mesh_15_8_io_in_last_1),
    .io_out_a_0(mesh_15_8_io_out_a_0),
    .io_out_a_1(mesh_15_8_io_out_a_1),
    .io_out_c_0(mesh_15_8_io_out_c_0),
    .io_out_c_1(mesh_15_8_io_out_c_1),
    .io_out_b_0(mesh_15_8_io_out_b_0),
    .io_out_b_1(mesh_15_8_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_8_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_8_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_8_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_8_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_8_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_8_io_out_control_1_shift),
    .io_out_id_0(mesh_15_8_io_out_id_0),
    .io_out_id_1(mesh_15_8_io_out_id_1),
    .io_out_last_0(mesh_15_8_io_out_last_0),
    .io_out_last_1(mesh_15_8_io_out_last_1),
    .io_in_valid_0(mesh_15_8_io_in_valid_0),
    .io_in_valid_1(mesh_15_8_io_in_valid_1),
    .io_out_valid_0(mesh_15_8_io_out_valid_0),
    .io_out_valid_1(mesh_15_8_io_out_valid_1)
  );
  Tile_240 mesh_15_9 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_9_clock),
    .io_in_a_0(mesh_15_9_io_in_a_0),
    .io_in_a_1(mesh_15_9_io_in_a_1),
    .io_in_b_0(mesh_15_9_io_in_b_0),
    .io_in_b_1(mesh_15_9_io_in_b_1),
    .io_in_d_0(mesh_15_9_io_in_d_0),
    .io_in_d_1(mesh_15_9_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_9_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_9_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_9_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_9_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_9_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_9_io_in_control_1_shift),
    .io_in_id_0(mesh_15_9_io_in_id_0),
    .io_in_id_1(mesh_15_9_io_in_id_1),
    .io_in_last_0(mesh_15_9_io_in_last_0),
    .io_in_last_1(mesh_15_9_io_in_last_1),
    .io_out_a_0(mesh_15_9_io_out_a_0),
    .io_out_a_1(mesh_15_9_io_out_a_1),
    .io_out_c_0(mesh_15_9_io_out_c_0),
    .io_out_c_1(mesh_15_9_io_out_c_1),
    .io_out_b_0(mesh_15_9_io_out_b_0),
    .io_out_b_1(mesh_15_9_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_9_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_9_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_9_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_9_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_9_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_9_io_out_control_1_shift),
    .io_out_id_0(mesh_15_9_io_out_id_0),
    .io_out_id_1(mesh_15_9_io_out_id_1),
    .io_out_last_0(mesh_15_9_io_out_last_0),
    .io_out_last_1(mesh_15_9_io_out_last_1),
    .io_in_valid_0(mesh_15_9_io_in_valid_0),
    .io_in_valid_1(mesh_15_9_io_in_valid_1),
    .io_out_valid_0(mesh_15_9_io_out_valid_0),
    .io_out_valid_1(mesh_15_9_io_out_valid_1)
  );
  Tile_240 mesh_15_10 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_10_clock),
    .io_in_a_0(mesh_15_10_io_in_a_0),
    .io_in_a_1(mesh_15_10_io_in_a_1),
    .io_in_b_0(mesh_15_10_io_in_b_0),
    .io_in_b_1(mesh_15_10_io_in_b_1),
    .io_in_d_0(mesh_15_10_io_in_d_0),
    .io_in_d_1(mesh_15_10_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_10_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_10_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_10_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_10_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_10_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_10_io_in_control_1_shift),
    .io_in_id_0(mesh_15_10_io_in_id_0),
    .io_in_id_1(mesh_15_10_io_in_id_1),
    .io_in_last_0(mesh_15_10_io_in_last_0),
    .io_in_last_1(mesh_15_10_io_in_last_1),
    .io_out_a_0(mesh_15_10_io_out_a_0),
    .io_out_a_1(mesh_15_10_io_out_a_1),
    .io_out_c_0(mesh_15_10_io_out_c_0),
    .io_out_c_1(mesh_15_10_io_out_c_1),
    .io_out_b_0(mesh_15_10_io_out_b_0),
    .io_out_b_1(mesh_15_10_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_10_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_10_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_10_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_10_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_10_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_10_io_out_control_1_shift),
    .io_out_id_0(mesh_15_10_io_out_id_0),
    .io_out_id_1(mesh_15_10_io_out_id_1),
    .io_out_last_0(mesh_15_10_io_out_last_0),
    .io_out_last_1(mesh_15_10_io_out_last_1),
    .io_in_valid_0(mesh_15_10_io_in_valid_0),
    .io_in_valid_1(mesh_15_10_io_in_valid_1),
    .io_out_valid_0(mesh_15_10_io_out_valid_0),
    .io_out_valid_1(mesh_15_10_io_out_valid_1)
  );
  Tile_240 mesh_15_11 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_11_clock),
    .io_in_a_0(mesh_15_11_io_in_a_0),
    .io_in_a_1(mesh_15_11_io_in_a_1),
    .io_in_b_0(mesh_15_11_io_in_b_0),
    .io_in_b_1(mesh_15_11_io_in_b_1),
    .io_in_d_0(mesh_15_11_io_in_d_0),
    .io_in_d_1(mesh_15_11_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_11_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_11_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_11_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_11_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_11_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_11_io_in_control_1_shift),
    .io_in_id_0(mesh_15_11_io_in_id_0),
    .io_in_id_1(mesh_15_11_io_in_id_1),
    .io_in_last_0(mesh_15_11_io_in_last_0),
    .io_in_last_1(mesh_15_11_io_in_last_1),
    .io_out_a_0(mesh_15_11_io_out_a_0),
    .io_out_a_1(mesh_15_11_io_out_a_1),
    .io_out_c_0(mesh_15_11_io_out_c_0),
    .io_out_c_1(mesh_15_11_io_out_c_1),
    .io_out_b_0(mesh_15_11_io_out_b_0),
    .io_out_b_1(mesh_15_11_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_11_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_11_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_11_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_11_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_11_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_11_io_out_control_1_shift),
    .io_out_id_0(mesh_15_11_io_out_id_0),
    .io_out_id_1(mesh_15_11_io_out_id_1),
    .io_out_last_0(mesh_15_11_io_out_last_0),
    .io_out_last_1(mesh_15_11_io_out_last_1),
    .io_in_valid_0(mesh_15_11_io_in_valid_0),
    .io_in_valid_1(mesh_15_11_io_in_valid_1),
    .io_out_valid_0(mesh_15_11_io_out_valid_0),
    .io_out_valid_1(mesh_15_11_io_out_valid_1)
  );
  Tile_240 mesh_15_12 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_12_clock),
    .io_in_a_0(mesh_15_12_io_in_a_0),
    .io_in_a_1(mesh_15_12_io_in_a_1),
    .io_in_b_0(mesh_15_12_io_in_b_0),
    .io_in_b_1(mesh_15_12_io_in_b_1),
    .io_in_d_0(mesh_15_12_io_in_d_0),
    .io_in_d_1(mesh_15_12_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_12_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_12_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_12_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_12_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_12_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_12_io_in_control_1_shift),
    .io_in_id_0(mesh_15_12_io_in_id_0),
    .io_in_id_1(mesh_15_12_io_in_id_1),
    .io_in_last_0(mesh_15_12_io_in_last_0),
    .io_in_last_1(mesh_15_12_io_in_last_1),
    .io_out_a_0(mesh_15_12_io_out_a_0),
    .io_out_a_1(mesh_15_12_io_out_a_1),
    .io_out_c_0(mesh_15_12_io_out_c_0),
    .io_out_c_1(mesh_15_12_io_out_c_1),
    .io_out_b_0(mesh_15_12_io_out_b_0),
    .io_out_b_1(mesh_15_12_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_12_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_12_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_12_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_12_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_12_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_12_io_out_control_1_shift),
    .io_out_id_0(mesh_15_12_io_out_id_0),
    .io_out_id_1(mesh_15_12_io_out_id_1),
    .io_out_last_0(mesh_15_12_io_out_last_0),
    .io_out_last_1(mesh_15_12_io_out_last_1),
    .io_in_valid_0(mesh_15_12_io_in_valid_0),
    .io_in_valid_1(mesh_15_12_io_in_valid_1),
    .io_out_valid_0(mesh_15_12_io_out_valid_0),
    .io_out_valid_1(mesh_15_12_io_out_valid_1)
  );
  Tile_240 mesh_15_13 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_13_clock),
    .io_in_a_0(mesh_15_13_io_in_a_0),
    .io_in_a_1(mesh_15_13_io_in_a_1),
    .io_in_b_0(mesh_15_13_io_in_b_0),
    .io_in_b_1(mesh_15_13_io_in_b_1),
    .io_in_d_0(mesh_15_13_io_in_d_0),
    .io_in_d_1(mesh_15_13_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_13_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_13_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_13_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_13_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_13_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_13_io_in_control_1_shift),
    .io_in_id_0(mesh_15_13_io_in_id_0),
    .io_in_id_1(mesh_15_13_io_in_id_1),
    .io_in_last_0(mesh_15_13_io_in_last_0),
    .io_in_last_1(mesh_15_13_io_in_last_1),
    .io_out_a_0(mesh_15_13_io_out_a_0),
    .io_out_a_1(mesh_15_13_io_out_a_1),
    .io_out_c_0(mesh_15_13_io_out_c_0),
    .io_out_c_1(mesh_15_13_io_out_c_1),
    .io_out_b_0(mesh_15_13_io_out_b_0),
    .io_out_b_1(mesh_15_13_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_13_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_13_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_13_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_13_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_13_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_13_io_out_control_1_shift),
    .io_out_id_0(mesh_15_13_io_out_id_0),
    .io_out_id_1(mesh_15_13_io_out_id_1),
    .io_out_last_0(mesh_15_13_io_out_last_0),
    .io_out_last_1(mesh_15_13_io_out_last_1),
    .io_in_valid_0(mesh_15_13_io_in_valid_0),
    .io_in_valid_1(mesh_15_13_io_in_valid_1),
    .io_out_valid_0(mesh_15_13_io_out_valid_0),
    .io_out_valid_1(mesh_15_13_io_out_valid_1)
  );
  Tile_240 mesh_15_14 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_14_clock),
    .io_in_a_0(mesh_15_14_io_in_a_0),
    .io_in_a_1(mesh_15_14_io_in_a_1),
    .io_in_b_0(mesh_15_14_io_in_b_0),
    .io_in_b_1(mesh_15_14_io_in_b_1),
    .io_in_d_0(mesh_15_14_io_in_d_0),
    .io_in_d_1(mesh_15_14_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_14_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_14_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_14_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_14_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_14_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_14_io_in_control_1_shift),
    .io_in_id_0(mesh_15_14_io_in_id_0),
    .io_in_id_1(mesh_15_14_io_in_id_1),
    .io_in_last_0(mesh_15_14_io_in_last_0),
    .io_in_last_1(mesh_15_14_io_in_last_1),
    .io_out_a_0(mesh_15_14_io_out_a_0),
    .io_out_a_1(mesh_15_14_io_out_a_1),
    .io_out_c_0(mesh_15_14_io_out_c_0),
    .io_out_c_1(mesh_15_14_io_out_c_1),
    .io_out_b_0(mesh_15_14_io_out_b_0),
    .io_out_b_1(mesh_15_14_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_14_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_14_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_14_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_14_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_14_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_14_io_out_control_1_shift),
    .io_out_id_0(mesh_15_14_io_out_id_0),
    .io_out_id_1(mesh_15_14_io_out_id_1),
    .io_out_last_0(mesh_15_14_io_out_last_0),
    .io_out_last_1(mesh_15_14_io_out_last_1),
    .io_in_valid_0(mesh_15_14_io_in_valid_0),
    .io_in_valid_1(mesh_15_14_io_in_valid_1),
    .io_out_valid_0(mesh_15_14_io_out_valid_0),
    .io_out_valid_1(mesh_15_14_io_out_valid_1)
  );
  Tile_240 mesh_15_15 ( // @[src/main/scala/gemmini/Mesh.scala 39:71]
    .clock(mesh_15_15_clock),
    .io_in_a_0(mesh_15_15_io_in_a_0),
    .io_in_a_1(mesh_15_15_io_in_a_1),
    .io_in_b_0(mesh_15_15_io_in_b_0),
    .io_in_b_1(mesh_15_15_io_in_b_1),
    .io_in_d_0(mesh_15_15_io_in_d_0),
    .io_in_d_1(mesh_15_15_io_in_d_1),
    .io_in_control_0_dataflow(mesh_15_15_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_15_15_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_15_15_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_15_15_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_15_15_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_15_15_io_in_control_1_shift),
    .io_in_id_0(mesh_15_15_io_in_id_0),
    .io_in_id_1(mesh_15_15_io_in_id_1),
    .io_in_last_0(mesh_15_15_io_in_last_0),
    .io_in_last_1(mesh_15_15_io_in_last_1),
    .io_out_a_0(mesh_15_15_io_out_a_0),
    .io_out_a_1(mesh_15_15_io_out_a_1),
    .io_out_c_0(mesh_15_15_io_out_c_0),
    .io_out_c_1(mesh_15_15_io_out_c_1),
    .io_out_b_0(mesh_15_15_io_out_b_0),
    .io_out_b_1(mesh_15_15_io_out_b_1),
    .io_out_control_0_dataflow(mesh_15_15_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_15_15_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_15_15_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_15_15_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_15_15_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_15_15_io_out_control_1_shift),
    .io_out_id_0(mesh_15_15_io_out_id_0),
    .io_out_id_1(mesh_15_15_io_out_id_1),
    .io_out_last_0(mesh_15_15_io_out_last_0),
    .io_out_last_1(mesh_15_15_io_out_last_1),
    .io_in_valid_0(mesh_15_15_io_in_valid_0),
    .io_in_valid_1(mesh_15_15_io_in_valid_1),
    .io_out_valid_0(mesh_15_15_io_out_valid_0),
    .io_out_valid_1(mesh_15_15_io_out_valid_1)
  );
  assign io_out_b_0_0 = mesh_15_0_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_0_1 = mesh_15_0_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_1_0 = mesh_15_1_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_1_1 = mesh_15_1_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_2_0 = mesh_15_2_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_2_1 = mesh_15_2_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_3_0 = mesh_15_3_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_3_1 = mesh_15_3_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_4_0 = mesh_15_4_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_4_1 = mesh_15_4_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_5_0 = mesh_15_5_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_5_1 = mesh_15_5_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_6_0 = mesh_15_6_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_6_1 = mesh_15_6_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_7_0 = mesh_15_7_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_7_1 = mesh_15_7_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_8_0 = mesh_15_8_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_8_1 = mesh_15_8_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_9_0 = mesh_15_9_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_9_1 = mesh_15_9_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_10_0 = mesh_15_10_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_10_1 = mesh_15_10_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_11_0 = mesh_15_11_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_11_1 = mesh_15_11_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_12_0 = mesh_15_12_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_12_1 = mesh_15_12_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_13_0 = mesh_15_13_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_13_1 = mesh_15_13_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_14_0 = mesh_15_14_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_14_1 = mesh_15_14_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_15_0 = mesh_15_15_io_out_b_0; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_b_15_1 = mesh_15_15_io_out_b_1; // @[src/main/scala/gemmini/Mesh.scala 122:7]
  assign io_out_c_0_0 = mesh_15_0_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_0_1 = mesh_15_0_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_1_0 = mesh_15_1_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_1_1 = mesh_15_1_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_2_0 = mesh_15_2_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_2_1 = mesh_15_2_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_3_0 = mesh_15_3_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_3_1 = mesh_15_3_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_4_0 = mesh_15_4_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_4_1 = mesh_15_4_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_5_0 = mesh_15_5_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_5_1 = mesh_15_5_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_6_0 = mesh_15_6_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_6_1 = mesh_15_6_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_7_0 = mesh_15_7_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_7_1 = mesh_15_7_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_8_0 = mesh_15_8_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_8_1 = mesh_15_8_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_9_0 = mesh_15_9_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_9_1 = mesh_15_9_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_10_0 = mesh_15_10_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_10_1 = mesh_15_10_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_11_0 = mesh_15_11_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_11_1 = mesh_15_11_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_12_0 = mesh_15_12_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_12_1 = mesh_15_12_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_13_0 = mesh_15_13_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_13_1 = mesh_15_13_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_14_0 = mesh_15_14_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_14_1 = mesh_15_14_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_15_0 = mesh_15_15_io_out_c_0; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_c_15_1 = mesh_15_15_io_out_c_1; // @[src/main/scala/gemmini/Mesh.scala 123:7]
  assign io_out_valid_0_0 = mesh_15_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_0_1 = mesh_15_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_1_0 = mesh_15_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_1_1 = mesh_15_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_2_0 = mesh_15_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_2_1 = mesh_15_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_3_0 = mesh_15_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_3_1 = mesh_15_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_4_0 = mesh_15_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_4_1 = mesh_15_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_5_0 = mesh_15_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_5_1 = mesh_15_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_6_0 = mesh_15_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_6_1 = mesh_15_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_7_0 = mesh_15_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_7_1 = mesh_15_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_8_0 = mesh_15_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_8_1 = mesh_15_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_9_0 = mesh_15_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_9_1 = mesh_15_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_10_0 = mesh_15_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_10_1 = mesh_15_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_11_0 = mesh_15_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_11_1 = mesh_15_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_12_0 = mesh_15_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_12_1 = mesh_15_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_13_0 = mesh_15_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_13_1 = mesh_15_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_14_0 = mesh_15_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_14_1 = mesh_15_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_15_0 = mesh_15_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_valid_15_1 = mesh_15_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 124:7]
  assign io_out_control_0_0_dataflow = mesh_15_0_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_0_0_propagate = mesh_15_0_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_0_0_shift = mesh_15_0_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_0_1_dataflow = mesh_15_0_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_0_1_propagate = mesh_15_0_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_0_1_shift = mesh_15_0_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_1_0_dataflow = mesh_15_1_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_1_0_propagate = mesh_15_1_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_1_0_shift = mesh_15_1_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_1_1_dataflow = mesh_15_1_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_1_1_propagate = mesh_15_1_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_1_1_shift = mesh_15_1_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_2_0_dataflow = mesh_15_2_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_2_0_propagate = mesh_15_2_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_2_0_shift = mesh_15_2_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_2_1_dataflow = mesh_15_2_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_2_1_propagate = mesh_15_2_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_2_1_shift = mesh_15_2_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_3_0_dataflow = mesh_15_3_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_3_0_propagate = mesh_15_3_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_3_0_shift = mesh_15_3_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_3_1_dataflow = mesh_15_3_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_3_1_propagate = mesh_15_3_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_3_1_shift = mesh_15_3_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_4_0_dataflow = mesh_15_4_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_4_0_propagate = mesh_15_4_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_4_0_shift = mesh_15_4_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_4_1_dataflow = mesh_15_4_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_4_1_propagate = mesh_15_4_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_4_1_shift = mesh_15_4_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_5_0_dataflow = mesh_15_5_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_5_0_propagate = mesh_15_5_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_5_0_shift = mesh_15_5_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_5_1_dataflow = mesh_15_5_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_5_1_propagate = mesh_15_5_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_5_1_shift = mesh_15_5_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_6_0_dataflow = mesh_15_6_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_6_0_propagate = mesh_15_6_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_6_0_shift = mesh_15_6_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_6_1_dataflow = mesh_15_6_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_6_1_propagate = mesh_15_6_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_6_1_shift = mesh_15_6_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_7_0_dataflow = mesh_15_7_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_7_0_propagate = mesh_15_7_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_7_0_shift = mesh_15_7_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_7_1_dataflow = mesh_15_7_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_7_1_propagate = mesh_15_7_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_7_1_shift = mesh_15_7_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_8_0_dataflow = mesh_15_8_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_8_0_propagate = mesh_15_8_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_8_0_shift = mesh_15_8_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_8_1_dataflow = mesh_15_8_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_8_1_propagate = mesh_15_8_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_8_1_shift = mesh_15_8_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_9_0_dataflow = mesh_15_9_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_9_0_propagate = mesh_15_9_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_9_0_shift = mesh_15_9_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_9_1_dataflow = mesh_15_9_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_9_1_propagate = mesh_15_9_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_9_1_shift = mesh_15_9_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_10_0_dataflow = mesh_15_10_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_10_0_propagate = mesh_15_10_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_10_0_shift = mesh_15_10_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_10_1_dataflow = mesh_15_10_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_10_1_propagate = mesh_15_10_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_10_1_shift = mesh_15_10_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_11_0_dataflow = mesh_15_11_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_11_0_propagate = mesh_15_11_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_11_0_shift = mesh_15_11_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_11_1_dataflow = mesh_15_11_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_11_1_propagate = mesh_15_11_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_11_1_shift = mesh_15_11_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_12_0_dataflow = mesh_15_12_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_12_0_propagate = mesh_15_12_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_12_0_shift = mesh_15_12_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_12_1_dataflow = mesh_15_12_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_12_1_propagate = mesh_15_12_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_12_1_shift = mesh_15_12_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_13_0_dataflow = mesh_15_13_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_13_0_propagate = mesh_15_13_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_13_0_shift = mesh_15_13_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_13_1_dataflow = mesh_15_13_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_13_1_propagate = mesh_15_13_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_13_1_shift = mesh_15_13_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_14_0_dataflow = mesh_15_14_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_14_0_propagate = mesh_15_14_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_14_0_shift = mesh_15_14_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_14_1_dataflow = mesh_15_14_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_14_1_propagate = mesh_15_14_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_14_1_shift = mesh_15_14_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_15_0_dataflow = mesh_15_15_io_out_control_0_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_15_0_propagate = mesh_15_15_io_out_control_0_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_15_0_shift = mesh_15_15_io_out_control_0_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_15_1_dataflow = mesh_15_15_io_out_control_1_dataflow; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_15_1_propagate = mesh_15_15_io_out_control_1_propagate; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_control_15_1_shift = mesh_15_15_io_out_control_1_shift; // @[src/main/scala/gemmini/Mesh.scala 125:10]
  assign io_out_id_0_0 = mesh_15_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_0_1 = mesh_15_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_1_0 = mesh_15_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_1_1 = mesh_15_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_2_0 = mesh_15_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_2_1 = mesh_15_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_3_0 = mesh_15_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_3_1 = mesh_15_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_4_0 = mesh_15_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_4_1 = mesh_15_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_5_0 = mesh_15_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_5_1 = mesh_15_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_6_0 = mesh_15_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_6_1 = mesh_15_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_7_0 = mesh_15_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_7_1 = mesh_15_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_8_0 = mesh_15_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_8_1 = mesh_15_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_9_0 = mesh_15_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_9_1 = mesh_15_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_10_0 = mesh_15_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_10_1 = mesh_15_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_11_0 = mesh_15_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_11_1 = mesh_15_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_12_0 = mesh_15_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_12_1 = mesh_15_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_13_0 = mesh_15_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_13_1 = mesh_15_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_14_0 = mesh_15_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_14_1 = mesh_15_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_15_0 = mesh_15_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_id_15_1 = mesh_15_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 126:8]
  assign io_out_last_0_0 = mesh_15_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_0_1 = mesh_15_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_1_0 = mesh_15_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_1_1 = mesh_15_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_2_0 = mesh_15_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_2_1 = mesh_15_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_3_0 = mesh_15_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_3_1 = mesh_15_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_4_0 = mesh_15_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_4_1 = mesh_15_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_5_0 = mesh_15_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_5_1 = mesh_15_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_6_0 = mesh_15_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_6_1 = mesh_15_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_7_0 = mesh_15_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_7_1 = mesh_15_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_8_0 = mesh_15_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_8_1 = mesh_15_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_9_0 = mesh_15_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_9_1 = mesh_15_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_10_0 = mesh_15_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_10_1 = mesh_15_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_11_0 = mesh_15_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_11_1 = mesh_15_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_12_0 = mesh_15_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_12_1 = mesh_15_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_13_0 = mesh_15_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_13_1 = mesh_15_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_14_0 = mesh_15_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_14_1 = mesh_15_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_15_0 = mesh_15_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign io_out_last_15_1 = mesh_15_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 127:10]
  assign mesh_0_0_clock = clock;
  assign mesh_0_0_io_in_a_0 = r__0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_0_io_in_a_1 = r__1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_0_io_in_b_0 = {{12{pipe_b__0[7]}},pipe_b__0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_0_io_in_b_1 = {{12{pipe_b__1[7]}},pipe_b__1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_0_io_in_d_0 = {{12{pipe_b_256_0[7]}},pipe_b_256_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_0_io_in_d_1 = {{12{pipe_b_256_1[7]}},pipe_b_256_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_0_io_in_control_0_dataflow = mesh_0_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_0_io_in_control_0_propagate = mesh_0_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_0_io_in_control_0_shift = mesh_0_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_0_io_in_control_1_dataflow = mesh_0_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_0_io_in_control_1_propagate = mesh_0_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_0_io_in_control_1_shift = mesh_0_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_0_io_in_id_0 = r_512_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_0_io_in_id_1 = r_512_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_0_io_in_last_0 = r_768_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_0_io_in_last_1 = r_768_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_0_io_in_valid_0 = r_256_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_0_io_in_valid_1 = r_256_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_1_clock = clock;
  assign mesh_0_1_io_in_a_0 = r_1_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_1_io_in_a_1 = r_1_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_1_io_in_b_0 = {{12{pipe_b_16_0[7]}},pipe_b_16_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_1_io_in_b_1 = {{12{pipe_b_16_1[7]}},pipe_b_16_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_1_io_in_d_0 = {{12{pipe_b_272_0[7]}},pipe_b_272_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_1_io_in_d_1 = {{12{pipe_b_272_1[7]}},pipe_b_272_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_1_io_in_control_0_dataflow = mesh_0_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_1_io_in_control_0_propagate = mesh_0_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_1_io_in_control_0_shift = mesh_0_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_1_io_in_control_1_dataflow = mesh_0_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_1_io_in_control_1_propagate = mesh_0_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_1_io_in_control_1_shift = mesh_0_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_1_io_in_id_0 = r_528_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_1_io_in_id_1 = r_528_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_1_io_in_last_0 = r_784_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_1_io_in_last_1 = r_784_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_1_io_in_valid_0 = r_272_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_1_io_in_valid_1 = r_272_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_2_clock = clock;
  assign mesh_0_2_io_in_a_0 = r_2_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_2_io_in_a_1 = r_2_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_2_io_in_b_0 = {{12{pipe_b_32_0[7]}},pipe_b_32_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_2_io_in_b_1 = {{12{pipe_b_32_1[7]}},pipe_b_32_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_2_io_in_d_0 = {{12{pipe_b_288_0[7]}},pipe_b_288_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_2_io_in_d_1 = {{12{pipe_b_288_1[7]}},pipe_b_288_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_2_io_in_control_0_dataflow = mesh_0_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_2_io_in_control_0_propagate = mesh_0_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_2_io_in_control_0_shift = mesh_0_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_2_io_in_control_1_dataflow = mesh_0_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_2_io_in_control_1_propagate = mesh_0_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_2_io_in_control_1_shift = mesh_0_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_2_io_in_id_0 = r_544_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_2_io_in_id_1 = r_544_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_2_io_in_last_0 = r_800_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_2_io_in_last_1 = r_800_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_2_io_in_valid_0 = r_288_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_2_io_in_valid_1 = r_288_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_3_clock = clock;
  assign mesh_0_3_io_in_a_0 = r_3_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_3_io_in_a_1 = r_3_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_3_io_in_b_0 = {{12{pipe_b_48_0[7]}},pipe_b_48_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_3_io_in_b_1 = {{12{pipe_b_48_1[7]}},pipe_b_48_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_3_io_in_d_0 = {{12{pipe_b_304_0[7]}},pipe_b_304_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_3_io_in_d_1 = {{12{pipe_b_304_1[7]}},pipe_b_304_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_3_io_in_control_0_dataflow = mesh_0_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_3_io_in_control_0_propagate = mesh_0_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_3_io_in_control_0_shift = mesh_0_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_3_io_in_control_1_dataflow = mesh_0_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_3_io_in_control_1_propagate = mesh_0_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_3_io_in_control_1_shift = mesh_0_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_3_io_in_id_0 = r_560_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_3_io_in_id_1 = r_560_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_3_io_in_last_0 = r_816_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_3_io_in_last_1 = r_816_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_3_io_in_valid_0 = r_304_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_3_io_in_valid_1 = r_304_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_4_clock = clock;
  assign mesh_0_4_io_in_a_0 = r_4_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_4_io_in_a_1 = r_4_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_4_io_in_b_0 = {{12{pipe_b_64_0[7]}},pipe_b_64_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_4_io_in_b_1 = {{12{pipe_b_64_1[7]}},pipe_b_64_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_4_io_in_d_0 = {{12{pipe_b_320_0[7]}},pipe_b_320_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_4_io_in_d_1 = {{12{pipe_b_320_1[7]}},pipe_b_320_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_4_io_in_control_0_dataflow = mesh_0_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_4_io_in_control_0_propagate = mesh_0_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_4_io_in_control_0_shift = mesh_0_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_4_io_in_control_1_dataflow = mesh_0_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_4_io_in_control_1_propagate = mesh_0_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_4_io_in_control_1_shift = mesh_0_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_4_io_in_id_0 = r_576_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_4_io_in_id_1 = r_576_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_4_io_in_last_0 = r_832_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_4_io_in_last_1 = r_832_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_4_io_in_valid_0 = r_320_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_4_io_in_valid_1 = r_320_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_5_clock = clock;
  assign mesh_0_5_io_in_a_0 = r_5_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_5_io_in_a_1 = r_5_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_5_io_in_b_0 = {{12{pipe_b_80_0[7]}},pipe_b_80_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_5_io_in_b_1 = {{12{pipe_b_80_1[7]}},pipe_b_80_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_5_io_in_d_0 = {{12{pipe_b_336_0[7]}},pipe_b_336_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_5_io_in_d_1 = {{12{pipe_b_336_1[7]}},pipe_b_336_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_5_io_in_control_0_dataflow = mesh_0_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_5_io_in_control_0_propagate = mesh_0_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_5_io_in_control_0_shift = mesh_0_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_5_io_in_control_1_dataflow = mesh_0_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_5_io_in_control_1_propagate = mesh_0_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_5_io_in_control_1_shift = mesh_0_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_5_io_in_id_0 = r_592_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_5_io_in_id_1 = r_592_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_5_io_in_last_0 = r_848_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_5_io_in_last_1 = r_848_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_5_io_in_valid_0 = r_336_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_5_io_in_valid_1 = r_336_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_6_clock = clock;
  assign mesh_0_6_io_in_a_0 = r_6_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_6_io_in_a_1 = r_6_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_6_io_in_b_0 = {{12{pipe_b_96_0[7]}},pipe_b_96_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_6_io_in_b_1 = {{12{pipe_b_96_1[7]}},pipe_b_96_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_6_io_in_d_0 = {{12{pipe_b_352_0[7]}},pipe_b_352_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_6_io_in_d_1 = {{12{pipe_b_352_1[7]}},pipe_b_352_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_6_io_in_control_0_dataflow = mesh_0_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_6_io_in_control_0_propagate = mesh_0_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_6_io_in_control_0_shift = mesh_0_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_6_io_in_control_1_dataflow = mesh_0_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_6_io_in_control_1_propagate = mesh_0_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_6_io_in_control_1_shift = mesh_0_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_6_io_in_id_0 = r_608_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_6_io_in_id_1 = r_608_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_6_io_in_last_0 = r_864_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_6_io_in_last_1 = r_864_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_6_io_in_valid_0 = r_352_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_6_io_in_valid_1 = r_352_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_7_clock = clock;
  assign mesh_0_7_io_in_a_0 = r_7_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_7_io_in_a_1 = r_7_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_7_io_in_b_0 = {{12{pipe_b_112_0[7]}},pipe_b_112_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_7_io_in_b_1 = {{12{pipe_b_112_1[7]}},pipe_b_112_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_7_io_in_d_0 = {{12{pipe_b_368_0[7]}},pipe_b_368_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_7_io_in_d_1 = {{12{pipe_b_368_1[7]}},pipe_b_368_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_7_io_in_control_0_dataflow = mesh_0_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_7_io_in_control_0_propagate = mesh_0_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_7_io_in_control_0_shift = mesh_0_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_7_io_in_control_1_dataflow = mesh_0_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_7_io_in_control_1_propagate = mesh_0_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_7_io_in_control_1_shift = mesh_0_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_7_io_in_id_0 = r_624_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_7_io_in_id_1 = r_624_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_7_io_in_last_0 = r_880_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_7_io_in_last_1 = r_880_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_7_io_in_valid_0 = r_368_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_7_io_in_valid_1 = r_368_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_8_clock = clock;
  assign mesh_0_8_io_in_a_0 = r_8_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_8_io_in_a_1 = r_8_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_8_io_in_b_0 = {{12{pipe_b_128_0[7]}},pipe_b_128_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_8_io_in_b_1 = {{12{pipe_b_128_1[7]}},pipe_b_128_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_8_io_in_d_0 = {{12{pipe_b_384_0[7]}},pipe_b_384_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_8_io_in_d_1 = {{12{pipe_b_384_1[7]}},pipe_b_384_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_8_io_in_control_0_dataflow = mesh_0_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_8_io_in_control_0_propagate = mesh_0_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_8_io_in_control_0_shift = mesh_0_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_8_io_in_control_1_dataflow = mesh_0_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_8_io_in_control_1_propagate = mesh_0_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_8_io_in_control_1_shift = mesh_0_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_8_io_in_id_0 = r_640_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_8_io_in_id_1 = r_640_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_8_io_in_last_0 = r_896_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_8_io_in_last_1 = r_896_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_8_io_in_valid_0 = r_384_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_8_io_in_valid_1 = r_384_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_9_clock = clock;
  assign mesh_0_9_io_in_a_0 = r_9_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_9_io_in_a_1 = r_9_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_9_io_in_b_0 = {{12{pipe_b_144_0[7]}},pipe_b_144_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_9_io_in_b_1 = {{12{pipe_b_144_1[7]}},pipe_b_144_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_9_io_in_d_0 = {{12{pipe_b_400_0[7]}},pipe_b_400_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_9_io_in_d_1 = {{12{pipe_b_400_1[7]}},pipe_b_400_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_9_io_in_control_0_dataflow = mesh_0_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_9_io_in_control_0_propagate = mesh_0_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_9_io_in_control_0_shift = mesh_0_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_9_io_in_control_1_dataflow = mesh_0_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_9_io_in_control_1_propagate = mesh_0_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_9_io_in_control_1_shift = mesh_0_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_9_io_in_id_0 = r_656_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_9_io_in_id_1 = r_656_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_9_io_in_last_0 = r_912_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_9_io_in_last_1 = r_912_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_9_io_in_valid_0 = r_400_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_9_io_in_valid_1 = r_400_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_10_clock = clock;
  assign mesh_0_10_io_in_a_0 = r_10_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_10_io_in_a_1 = r_10_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_10_io_in_b_0 = {{12{pipe_b_160_0[7]}},pipe_b_160_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_10_io_in_b_1 = {{12{pipe_b_160_1[7]}},pipe_b_160_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_10_io_in_d_0 = {{12{pipe_b_416_0[7]}},pipe_b_416_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_10_io_in_d_1 = {{12{pipe_b_416_1[7]}},pipe_b_416_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_10_io_in_control_0_dataflow = mesh_0_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_10_io_in_control_0_propagate = mesh_0_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_10_io_in_control_0_shift = mesh_0_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_10_io_in_control_1_dataflow = mesh_0_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_10_io_in_control_1_propagate = mesh_0_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_10_io_in_control_1_shift = mesh_0_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_10_io_in_id_0 = r_672_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_10_io_in_id_1 = r_672_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_10_io_in_last_0 = r_928_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_10_io_in_last_1 = r_928_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_10_io_in_valid_0 = r_416_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_10_io_in_valid_1 = r_416_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_11_clock = clock;
  assign mesh_0_11_io_in_a_0 = r_11_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_11_io_in_a_1 = r_11_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_11_io_in_b_0 = {{12{pipe_b_176_0[7]}},pipe_b_176_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_11_io_in_b_1 = {{12{pipe_b_176_1[7]}},pipe_b_176_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_11_io_in_d_0 = {{12{pipe_b_432_0[7]}},pipe_b_432_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_11_io_in_d_1 = {{12{pipe_b_432_1[7]}},pipe_b_432_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_11_io_in_control_0_dataflow = mesh_0_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_11_io_in_control_0_propagate = mesh_0_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_11_io_in_control_0_shift = mesh_0_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_11_io_in_control_1_dataflow = mesh_0_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_11_io_in_control_1_propagate = mesh_0_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_11_io_in_control_1_shift = mesh_0_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_11_io_in_id_0 = r_688_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_11_io_in_id_1 = r_688_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_11_io_in_last_0 = r_944_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_11_io_in_last_1 = r_944_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_11_io_in_valid_0 = r_432_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_11_io_in_valid_1 = r_432_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_12_clock = clock;
  assign mesh_0_12_io_in_a_0 = r_12_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_12_io_in_a_1 = r_12_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_12_io_in_b_0 = {{12{pipe_b_192_0[7]}},pipe_b_192_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_12_io_in_b_1 = {{12{pipe_b_192_1[7]}},pipe_b_192_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_12_io_in_d_0 = {{12{pipe_b_448_0[7]}},pipe_b_448_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_12_io_in_d_1 = {{12{pipe_b_448_1[7]}},pipe_b_448_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_12_io_in_control_0_dataflow = mesh_0_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_12_io_in_control_0_propagate = mesh_0_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_12_io_in_control_0_shift = mesh_0_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_12_io_in_control_1_dataflow = mesh_0_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_12_io_in_control_1_propagate = mesh_0_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_12_io_in_control_1_shift = mesh_0_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_12_io_in_id_0 = r_704_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_12_io_in_id_1 = r_704_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_12_io_in_last_0 = r_960_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_12_io_in_last_1 = r_960_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_12_io_in_valid_0 = r_448_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_12_io_in_valid_1 = r_448_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_13_clock = clock;
  assign mesh_0_13_io_in_a_0 = r_13_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_13_io_in_a_1 = r_13_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_13_io_in_b_0 = {{12{pipe_b_208_0[7]}},pipe_b_208_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_13_io_in_b_1 = {{12{pipe_b_208_1[7]}},pipe_b_208_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_13_io_in_d_0 = {{12{pipe_b_464_0[7]}},pipe_b_464_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_13_io_in_d_1 = {{12{pipe_b_464_1[7]}},pipe_b_464_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_13_io_in_control_0_dataflow = mesh_0_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_13_io_in_control_0_propagate = mesh_0_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_13_io_in_control_0_shift = mesh_0_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_13_io_in_control_1_dataflow = mesh_0_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_13_io_in_control_1_propagate = mesh_0_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_13_io_in_control_1_shift = mesh_0_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_13_io_in_id_0 = r_720_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_13_io_in_id_1 = r_720_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_13_io_in_last_0 = r_976_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_13_io_in_last_1 = r_976_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_13_io_in_valid_0 = r_464_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_13_io_in_valid_1 = r_464_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_14_clock = clock;
  assign mesh_0_14_io_in_a_0 = r_14_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_14_io_in_a_1 = r_14_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_14_io_in_b_0 = {{12{pipe_b_224_0[7]}},pipe_b_224_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_14_io_in_b_1 = {{12{pipe_b_224_1[7]}},pipe_b_224_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_14_io_in_d_0 = {{12{pipe_b_480_0[7]}},pipe_b_480_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_14_io_in_d_1 = {{12{pipe_b_480_1[7]}},pipe_b_480_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_14_io_in_control_0_dataflow = mesh_0_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_14_io_in_control_0_propagate = mesh_0_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_14_io_in_control_0_shift = mesh_0_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_14_io_in_control_1_dataflow = mesh_0_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_14_io_in_control_1_propagate = mesh_0_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_14_io_in_control_1_shift = mesh_0_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_14_io_in_id_0 = r_736_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_14_io_in_id_1 = r_736_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_14_io_in_last_0 = r_992_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_14_io_in_last_1 = r_992_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_14_io_in_valid_0 = r_480_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_14_io_in_valid_1 = r_480_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_15_clock = clock;
  assign mesh_0_15_io_in_a_0 = r_15_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_15_io_in_a_1 = r_15_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_0_15_io_in_b_0 = {{12{pipe_b_240_0[7]}},pipe_b_240_0}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_15_io_in_b_1 = {{12{pipe_b_240_1[7]}},pipe_b_240_1}; // @[src/main/scala/gemmini/Mesh.scala 62:22]
  assign mesh_0_15_io_in_d_0 = {{12{pipe_b_496_0[7]}},pipe_b_496_0}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_15_io_in_d_1 = {{12{pipe_b_496_1[7]}},pipe_b_496_1}; // @[src/main/scala/gemmini/Mesh.scala 71:22]
  assign mesh_0_15_io_in_control_0_dataflow = mesh_0_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_15_io_in_control_0_propagate = mesh_0_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_15_io_in_control_0_shift = mesh_0_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_15_io_in_control_1_dataflow = mesh_0_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_15_io_in_control_1_propagate = mesh_0_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_15_io_in_control_1_shift = mesh_0_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_0_15_io_in_id_0 = r_752_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_15_io_in_id_1 = r_752_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_0_15_io_in_last_0 = r_1008_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_15_io_in_last_1 = r_1008_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_0_15_io_in_valid_0 = r_496_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_0_15_io_in_valid_1 = r_496_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_0_clock = clock;
  assign mesh_1_0_io_in_a_0 = r_16_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_0_io_in_a_1 = r_16_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_0_io_in_b_0 = pipe_b_1_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_b_1 = pipe_b_1_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_d_0 = pipe_b_257_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_d_1 = pipe_b_257_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_control_0_dataflow = mesh_1_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_control_0_propagate = mesh_1_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_control_0_shift = mesh_1_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_control_1_dataflow = mesh_1_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_control_1_propagate = mesh_1_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_control_1_shift = mesh_1_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_0_io_in_id_0 = r_513_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_0_io_in_id_1 = r_513_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_0_io_in_last_0 = r_769_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_0_io_in_last_1 = r_769_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_0_io_in_valid_0 = r_257_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_0_io_in_valid_1 = r_257_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_1_clock = clock;
  assign mesh_1_1_io_in_a_0 = r_17_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_1_io_in_a_1 = r_17_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_1_io_in_b_0 = pipe_b_17_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_b_1 = pipe_b_17_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_d_0 = pipe_b_273_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_d_1 = pipe_b_273_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_control_0_dataflow = mesh_1_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_control_0_propagate = mesh_1_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_control_0_shift = mesh_1_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_control_1_dataflow = mesh_1_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_control_1_propagate = mesh_1_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_control_1_shift = mesh_1_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_1_io_in_id_0 = r_529_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_1_io_in_id_1 = r_529_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_1_io_in_last_0 = r_785_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_1_io_in_last_1 = r_785_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_1_io_in_valid_0 = r_273_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_1_io_in_valid_1 = r_273_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_2_clock = clock;
  assign mesh_1_2_io_in_a_0 = r_18_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_2_io_in_a_1 = r_18_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_2_io_in_b_0 = pipe_b_33_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_b_1 = pipe_b_33_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_d_0 = pipe_b_289_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_d_1 = pipe_b_289_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_control_0_dataflow = mesh_1_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_control_0_propagate = mesh_1_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_control_0_shift = mesh_1_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_control_1_dataflow = mesh_1_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_control_1_propagate = mesh_1_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_control_1_shift = mesh_1_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_2_io_in_id_0 = r_545_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_2_io_in_id_1 = r_545_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_2_io_in_last_0 = r_801_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_2_io_in_last_1 = r_801_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_2_io_in_valid_0 = r_289_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_2_io_in_valid_1 = r_289_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_3_clock = clock;
  assign mesh_1_3_io_in_a_0 = r_19_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_3_io_in_a_1 = r_19_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_3_io_in_b_0 = pipe_b_49_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_b_1 = pipe_b_49_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_d_0 = pipe_b_305_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_d_1 = pipe_b_305_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_control_0_dataflow = mesh_1_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_control_0_propagate = mesh_1_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_control_0_shift = mesh_1_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_control_1_dataflow = mesh_1_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_control_1_propagate = mesh_1_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_control_1_shift = mesh_1_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_3_io_in_id_0 = r_561_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_3_io_in_id_1 = r_561_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_3_io_in_last_0 = r_817_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_3_io_in_last_1 = r_817_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_3_io_in_valid_0 = r_305_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_3_io_in_valid_1 = r_305_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_4_clock = clock;
  assign mesh_1_4_io_in_a_0 = r_20_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_4_io_in_a_1 = r_20_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_4_io_in_b_0 = pipe_b_65_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_b_1 = pipe_b_65_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_d_0 = pipe_b_321_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_d_1 = pipe_b_321_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_control_0_dataflow = mesh_1_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_control_0_propagate = mesh_1_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_control_0_shift = mesh_1_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_control_1_dataflow = mesh_1_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_control_1_propagate = mesh_1_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_control_1_shift = mesh_1_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_4_io_in_id_0 = r_577_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_4_io_in_id_1 = r_577_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_4_io_in_last_0 = r_833_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_4_io_in_last_1 = r_833_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_4_io_in_valid_0 = r_321_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_4_io_in_valid_1 = r_321_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_5_clock = clock;
  assign mesh_1_5_io_in_a_0 = r_21_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_5_io_in_a_1 = r_21_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_5_io_in_b_0 = pipe_b_81_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_b_1 = pipe_b_81_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_d_0 = pipe_b_337_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_d_1 = pipe_b_337_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_control_0_dataflow = mesh_1_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_control_0_propagate = mesh_1_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_control_0_shift = mesh_1_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_control_1_dataflow = mesh_1_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_control_1_propagate = mesh_1_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_control_1_shift = mesh_1_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_5_io_in_id_0 = r_593_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_5_io_in_id_1 = r_593_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_5_io_in_last_0 = r_849_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_5_io_in_last_1 = r_849_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_5_io_in_valid_0 = r_337_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_5_io_in_valid_1 = r_337_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_6_clock = clock;
  assign mesh_1_6_io_in_a_0 = r_22_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_6_io_in_a_1 = r_22_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_6_io_in_b_0 = pipe_b_97_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_b_1 = pipe_b_97_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_d_0 = pipe_b_353_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_d_1 = pipe_b_353_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_control_0_dataflow = mesh_1_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_control_0_propagate = mesh_1_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_control_0_shift = mesh_1_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_control_1_dataflow = mesh_1_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_control_1_propagate = mesh_1_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_control_1_shift = mesh_1_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_6_io_in_id_0 = r_609_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_6_io_in_id_1 = r_609_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_6_io_in_last_0 = r_865_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_6_io_in_last_1 = r_865_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_6_io_in_valid_0 = r_353_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_6_io_in_valid_1 = r_353_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_7_clock = clock;
  assign mesh_1_7_io_in_a_0 = r_23_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_7_io_in_a_1 = r_23_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_7_io_in_b_0 = pipe_b_113_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_b_1 = pipe_b_113_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_d_0 = pipe_b_369_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_d_1 = pipe_b_369_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_control_0_dataflow = mesh_1_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_control_0_propagate = mesh_1_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_control_0_shift = mesh_1_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_control_1_dataflow = mesh_1_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_control_1_propagate = mesh_1_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_control_1_shift = mesh_1_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_7_io_in_id_0 = r_625_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_7_io_in_id_1 = r_625_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_7_io_in_last_0 = r_881_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_7_io_in_last_1 = r_881_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_7_io_in_valid_0 = r_369_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_7_io_in_valid_1 = r_369_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_8_clock = clock;
  assign mesh_1_8_io_in_a_0 = r_24_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_8_io_in_a_1 = r_24_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_8_io_in_b_0 = pipe_b_129_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_b_1 = pipe_b_129_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_d_0 = pipe_b_385_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_d_1 = pipe_b_385_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_control_0_dataflow = mesh_1_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_control_0_propagate = mesh_1_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_control_0_shift = mesh_1_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_control_1_dataflow = mesh_1_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_control_1_propagate = mesh_1_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_control_1_shift = mesh_1_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_8_io_in_id_0 = r_641_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_8_io_in_id_1 = r_641_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_8_io_in_last_0 = r_897_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_8_io_in_last_1 = r_897_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_8_io_in_valid_0 = r_385_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_8_io_in_valid_1 = r_385_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_9_clock = clock;
  assign mesh_1_9_io_in_a_0 = r_25_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_9_io_in_a_1 = r_25_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_9_io_in_b_0 = pipe_b_145_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_b_1 = pipe_b_145_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_d_0 = pipe_b_401_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_d_1 = pipe_b_401_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_control_0_dataflow = mesh_1_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_control_0_propagate = mesh_1_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_control_0_shift = mesh_1_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_control_1_dataflow = mesh_1_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_control_1_propagate = mesh_1_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_control_1_shift = mesh_1_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_9_io_in_id_0 = r_657_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_9_io_in_id_1 = r_657_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_9_io_in_last_0 = r_913_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_9_io_in_last_1 = r_913_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_9_io_in_valid_0 = r_401_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_9_io_in_valid_1 = r_401_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_10_clock = clock;
  assign mesh_1_10_io_in_a_0 = r_26_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_10_io_in_a_1 = r_26_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_10_io_in_b_0 = pipe_b_161_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_b_1 = pipe_b_161_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_d_0 = pipe_b_417_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_d_1 = pipe_b_417_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_control_0_dataflow = mesh_1_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_control_0_propagate = mesh_1_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_control_0_shift = mesh_1_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_control_1_dataflow = mesh_1_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_control_1_propagate = mesh_1_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_control_1_shift = mesh_1_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_10_io_in_id_0 = r_673_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_10_io_in_id_1 = r_673_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_10_io_in_last_0 = r_929_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_10_io_in_last_1 = r_929_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_10_io_in_valid_0 = r_417_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_10_io_in_valid_1 = r_417_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_11_clock = clock;
  assign mesh_1_11_io_in_a_0 = r_27_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_11_io_in_a_1 = r_27_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_11_io_in_b_0 = pipe_b_177_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_b_1 = pipe_b_177_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_d_0 = pipe_b_433_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_d_1 = pipe_b_433_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_control_0_dataflow = mesh_1_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_control_0_propagate = mesh_1_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_control_0_shift = mesh_1_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_control_1_dataflow = mesh_1_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_control_1_propagate = mesh_1_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_control_1_shift = mesh_1_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_11_io_in_id_0 = r_689_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_11_io_in_id_1 = r_689_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_11_io_in_last_0 = r_945_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_11_io_in_last_1 = r_945_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_11_io_in_valid_0 = r_433_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_11_io_in_valid_1 = r_433_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_12_clock = clock;
  assign mesh_1_12_io_in_a_0 = r_28_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_12_io_in_a_1 = r_28_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_12_io_in_b_0 = pipe_b_193_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_b_1 = pipe_b_193_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_d_0 = pipe_b_449_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_d_1 = pipe_b_449_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_control_0_dataflow = mesh_1_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_control_0_propagate = mesh_1_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_control_0_shift = mesh_1_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_control_1_dataflow = mesh_1_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_control_1_propagate = mesh_1_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_control_1_shift = mesh_1_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_12_io_in_id_0 = r_705_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_12_io_in_id_1 = r_705_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_12_io_in_last_0 = r_961_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_12_io_in_last_1 = r_961_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_12_io_in_valid_0 = r_449_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_12_io_in_valid_1 = r_449_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_13_clock = clock;
  assign mesh_1_13_io_in_a_0 = r_29_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_13_io_in_a_1 = r_29_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_13_io_in_b_0 = pipe_b_209_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_b_1 = pipe_b_209_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_d_0 = pipe_b_465_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_d_1 = pipe_b_465_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_control_0_dataflow = mesh_1_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_control_0_propagate = mesh_1_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_control_0_shift = mesh_1_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_control_1_dataflow = mesh_1_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_control_1_propagate = mesh_1_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_control_1_shift = mesh_1_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_13_io_in_id_0 = r_721_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_13_io_in_id_1 = r_721_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_13_io_in_last_0 = r_977_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_13_io_in_last_1 = r_977_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_13_io_in_valid_0 = r_465_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_13_io_in_valid_1 = r_465_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_14_clock = clock;
  assign mesh_1_14_io_in_a_0 = r_30_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_14_io_in_a_1 = r_30_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_14_io_in_b_0 = pipe_b_225_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_b_1 = pipe_b_225_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_d_0 = pipe_b_481_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_d_1 = pipe_b_481_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_control_0_dataflow = mesh_1_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_control_0_propagate = mesh_1_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_control_0_shift = mesh_1_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_control_1_dataflow = mesh_1_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_control_1_propagate = mesh_1_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_control_1_shift = mesh_1_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_14_io_in_id_0 = r_737_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_14_io_in_id_1 = r_737_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_14_io_in_last_0 = r_993_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_14_io_in_last_1 = r_993_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_14_io_in_valid_0 = r_481_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_14_io_in_valid_1 = r_481_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_15_clock = clock;
  assign mesh_1_15_io_in_a_0 = r_31_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_15_io_in_a_1 = r_31_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_1_15_io_in_b_0 = pipe_b_241_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_b_1 = pipe_b_241_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_d_0 = pipe_b_497_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_d_1 = pipe_b_497_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_control_0_dataflow = mesh_1_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_control_0_propagate = mesh_1_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_control_0_shift = mesh_1_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_control_1_dataflow = mesh_1_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_control_1_propagate = mesh_1_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_control_1_shift = mesh_1_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_1_15_io_in_id_0 = r_753_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_15_io_in_id_1 = r_753_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_1_15_io_in_last_0 = r_1009_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_15_io_in_last_1 = r_1009_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_1_15_io_in_valid_0 = r_497_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_1_15_io_in_valid_1 = r_497_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_0_clock = clock;
  assign mesh_2_0_io_in_a_0 = r_32_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_0_io_in_a_1 = r_32_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_0_io_in_b_0 = pipe_b_2_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_b_1 = pipe_b_2_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_d_0 = pipe_b_258_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_d_1 = pipe_b_258_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_control_0_dataflow = mesh_2_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_control_0_propagate = mesh_2_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_control_0_shift = mesh_2_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_control_1_dataflow = mesh_2_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_control_1_propagate = mesh_2_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_control_1_shift = mesh_2_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_0_io_in_id_0 = r_514_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_0_io_in_id_1 = r_514_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_0_io_in_last_0 = r_770_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_0_io_in_last_1 = r_770_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_0_io_in_valid_0 = r_258_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_0_io_in_valid_1 = r_258_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_1_clock = clock;
  assign mesh_2_1_io_in_a_0 = r_33_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_1_io_in_a_1 = r_33_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_1_io_in_b_0 = pipe_b_18_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_b_1 = pipe_b_18_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_d_0 = pipe_b_274_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_d_1 = pipe_b_274_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_control_0_dataflow = mesh_2_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_control_0_propagate = mesh_2_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_control_0_shift = mesh_2_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_control_1_dataflow = mesh_2_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_control_1_propagate = mesh_2_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_control_1_shift = mesh_2_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_1_io_in_id_0 = r_530_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_1_io_in_id_1 = r_530_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_1_io_in_last_0 = r_786_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_1_io_in_last_1 = r_786_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_1_io_in_valid_0 = r_274_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_1_io_in_valid_1 = r_274_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_2_clock = clock;
  assign mesh_2_2_io_in_a_0 = r_34_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_2_io_in_a_1 = r_34_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_2_io_in_b_0 = pipe_b_34_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_b_1 = pipe_b_34_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_d_0 = pipe_b_290_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_d_1 = pipe_b_290_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_control_0_dataflow = mesh_2_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_control_0_propagate = mesh_2_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_control_0_shift = mesh_2_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_control_1_dataflow = mesh_2_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_control_1_propagate = mesh_2_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_control_1_shift = mesh_2_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_2_io_in_id_0 = r_546_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_2_io_in_id_1 = r_546_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_2_io_in_last_0 = r_802_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_2_io_in_last_1 = r_802_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_2_io_in_valid_0 = r_290_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_2_io_in_valid_1 = r_290_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_3_clock = clock;
  assign mesh_2_3_io_in_a_0 = r_35_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_3_io_in_a_1 = r_35_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_3_io_in_b_0 = pipe_b_50_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_b_1 = pipe_b_50_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_d_0 = pipe_b_306_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_d_1 = pipe_b_306_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_control_0_dataflow = mesh_2_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_control_0_propagate = mesh_2_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_control_0_shift = mesh_2_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_control_1_dataflow = mesh_2_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_control_1_propagate = mesh_2_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_control_1_shift = mesh_2_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_3_io_in_id_0 = r_562_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_3_io_in_id_1 = r_562_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_3_io_in_last_0 = r_818_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_3_io_in_last_1 = r_818_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_3_io_in_valid_0 = r_306_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_3_io_in_valid_1 = r_306_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_4_clock = clock;
  assign mesh_2_4_io_in_a_0 = r_36_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_4_io_in_a_1 = r_36_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_4_io_in_b_0 = pipe_b_66_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_b_1 = pipe_b_66_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_d_0 = pipe_b_322_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_d_1 = pipe_b_322_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_control_0_dataflow = mesh_2_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_control_0_propagate = mesh_2_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_control_0_shift = mesh_2_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_control_1_dataflow = mesh_2_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_control_1_propagate = mesh_2_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_control_1_shift = mesh_2_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_4_io_in_id_0 = r_578_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_4_io_in_id_1 = r_578_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_4_io_in_last_0 = r_834_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_4_io_in_last_1 = r_834_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_4_io_in_valid_0 = r_322_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_4_io_in_valid_1 = r_322_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_5_clock = clock;
  assign mesh_2_5_io_in_a_0 = r_37_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_5_io_in_a_1 = r_37_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_5_io_in_b_0 = pipe_b_82_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_b_1 = pipe_b_82_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_d_0 = pipe_b_338_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_d_1 = pipe_b_338_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_control_0_dataflow = mesh_2_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_control_0_propagate = mesh_2_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_control_0_shift = mesh_2_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_control_1_dataflow = mesh_2_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_control_1_propagate = mesh_2_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_control_1_shift = mesh_2_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_5_io_in_id_0 = r_594_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_5_io_in_id_1 = r_594_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_5_io_in_last_0 = r_850_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_5_io_in_last_1 = r_850_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_5_io_in_valid_0 = r_338_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_5_io_in_valid_1 = r_338_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_6_clock = clock;
  assign mesh_2_6_io_in_a_0 = r_38_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_6_io_in_a_1 = r_38_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_6_io_in_b_0 = pipe_b_98_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_b_1 = pipe_b_98_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_d_0 = pipe_b_354_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_d_1 = pipe_b_354_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_control_0_dataflow = mesh_2_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_control_0_propagate = mesh_2_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_control_0_shift = mesh_2_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_control_1_dataflow = mesh_2_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_control_1_propagate = mesh_2_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_control_1_shift = mesh_2_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_6_io_in_id_0 = r_610_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_6_io_in_id_1 = r_610_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_6_io_in_last_0 = r_866_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_6_io_in_last_1 = r_866_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_6_io_in_valid_0 = r_354_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_6_io_in_valid_1 = r_354_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_7_clock = clock;
  assign mesh_2_7_io_in_a_0 = r_39_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_7_io_in_a_1 = r_39_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_7_io_in_b_0 = pipe_b_114_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_b_1 = pipe_b_114_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_d_0 = pipe_b_370_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_d_1 = pipe_b_370_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_control_0_dataflow = mesh_2_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_control_0_propagate = mesh_2_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_control_0_shift = mesh_2_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_control_1_dataflow = mesh_2_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_control_1_propagate = mesh_2_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_control_1_shift = mesh_2_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_7_io_in_id_0 = r_626_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_7_io_in_id_1 = r_626_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_7_io_in_last_0 = r_882_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_7_io_in_last_1 = r_882_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_7_io_in_valid_0 = r_370_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_7_io_in_valid_1 = r_370_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_8_clock = clock;
  assign mesh_2_8_io_in_a_0 = r_40_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_8_io_in_a_1 = r_40_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_8_io_in_b_0 = pipe_b_130_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_b_1 = pipe_b_130_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_d_0 = pipe_b_386_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_d_1 = pipe_b_386_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_control_0_dataflow = mesh_2_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_control_0_propagate = mesh_2_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_control_0_shift = mesh_2_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_control_1_dataflow = mesh_2_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_control_1_propagate = mesh_2_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_control_1_shift = mesh_2_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_8_io_in_id_0 = r_642_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_8_io_in_id_1 = r_642_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_8_io_in_last_0 = r_898_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_8_io_in_last_1 = r_898_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_8_io_in_valid_0 = r_386_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_8_io_in_valid_1 = r_386_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_9_clock = clock;
  assign mesh_2_9_io_in_a_0 = r_41_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_9_io_in_a_1 = r_41_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_9_io_in_b_0 = pipe_b_146_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_b_1 = pipe_b_146_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_d_0 = pipe_b_402_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_d_1 = pipe_b_402_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_control_0_dataflow = mesh_2_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_control_0_propagate = mesh_2_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_control_0_shift = mesh_2_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_control_1_dataflow = mesh_2_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_control_1_propagate = mesh_2_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_control_1_shift = mesh_2_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_9_io_in_id_0 = r_658_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_9_io_in_id_1 = r_658_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_9_io_in_last_0 = r_914_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_9_io_in_last_1 = r_914_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_9_io_in_valid_0 = r_402_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_9_io_in_valid_1 = r_402_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_10_clock = clock;
  assign mesh_2_10_io_in_a_0 = r_42_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_10_io_in_a_1 = r_42_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_10_io_in_b_0 = pipe_b_162_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_b_1 = pipe_b_162_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_d_0 = pipe_b_418_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_d_1 = pipe_b_418_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_control_0_dataflow = mesh_2_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_control_0_propagate = mesh_2_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_control_0_shift = mesh_2_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_control_1_dataflow = mesh_2_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_control_1_propagate = mesh_2_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_control_1_shift = mesh_2_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_10_io_in_id_0 = r_674_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_10_io_in_id_1 = r_674_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_10_io_in_last_0 = r_930_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_10_io_in_last_1 = r_930_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_10_io_in_valid_0 = r_418_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_10_io_in_valid_1 = r_418_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_11_clock = clock;
  assign mesh_2_11_io_in_a_0 = r_43_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_11_io_in_a_1 = r_43_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_11_io_in_b_0 = pipe_b_178_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_b_1 = pipe_b_178_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_d_0 = pipe_b_434_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_d_1 = pipe_b_434_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_control_0_dataflow = mesh_2_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_control_0_propagate = mesh_2_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_control_0_shift = mesh_2_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_control_1_dataflow = mesh_2_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_control_1_propagate = mesh_2_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_control_1_shift = mesh_2_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_11_io_in_id_0 = r_690_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_11_io_in_id_1 = r_690_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_11_io_in_last_0 = r_946_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_11_io_in_last_1 = r_946_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_11_io_in_valid_0 = r_434_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_11_io_in_valid_1 = r_434_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_12_clock = clock;
  assign mesh_2_12_io_in_a_0 = r_44_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_12_io_in_a_1 = r_44_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_12_io_in_b_0 = pipe_b_194_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_b_1 = pipe_b_194_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_d_0 = pipe_b_450_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_d_1 = pipe_b_450_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_control_0_dataflow = mesh_2_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_control_0_propagate = mesh_2_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_control_0_shift = mesh_2_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_control_1_dataflow = mesh_2_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_control_1_propagate = mesh_2_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_control_1_shift = mesh_2_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_12_io_in_id_0 = r_706_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_12_io_in_id_1 = r_706_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_12_io_in_last_0 = r_962_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_12_io_in_last_1 = r_962_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_12_io_in_valid_0 = r_450_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_12_io_in_valid_1 = r_450_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_13_clock = clock;
  assign mesh_2_13_io_in_a_0 = r_45_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_13_io_in_a_1 = r_45_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_13_io_in_b_0 = pipe_b_210_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_b_1 = pipe_b_210_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_d_0 = pipe_b_466_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_d_1 = pipe_b_466_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_control_0_dataflow = mesh_2_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_control_0_propagate = mesh_2_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_control_0_shift = mesh_2_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_control_1_dataflow = mesh_2_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_control_1_propagate = mesh_2_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_control_1_shift = mesh_2_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_13_io_in_id_0 = r_722_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_13_io_in_id_1 = r_722_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_13_io_in_last_0 = r_978_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_13_io_in_last_1 = r_978_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_13_io_in_valid_0 = r_466_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_13_io_in_valid_1 = r_466_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_14_clock = clock;
  assign mesh_2_14_io_in_a_0 = r_46_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_14_io_in_a_1 = r_46_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_14_io_in_b_0 = pipe_b_226_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_b_1 = pipe_b_226_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_d_0 = pipe_b_482_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_d_1 = pipe_b_482_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_control_0_dataflow = mesh_2_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_control_0_propagate = mesh_2_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_control_0_shift = mesh_2_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_control_1_dataflow = mesh_2_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_control_1_propagate = mesh_2_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_control_1_shift = mesh_2_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_14_io_in_id_0 = r_738_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_14_io_in_id_1 = r_738_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_14_io_in_last_0 = r_994_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_14_io_in_last_1 = r_994_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_14_io_in_valid_0 = r_482_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_14_io_in_valid_1 = r_482_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_15_clock = clock;
  assign mesh_2_15_io_in_a_0 = r_47_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_15_io_in_a_1 = r_47_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_2_15_io_in_b_0 = pipe_b_242_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_b_1 = pipe_b_242_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_d_0 = pipe_b_498_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_d_1 = pipe_b_498_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_control_0_dataflow = mesh_2_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_control_0_propagate = mesh_2_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_control_0_shift = mesh_2_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_control_1_dataflow = mesh_2_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_control_1_propagate = mesh_2_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_control_1_shift = mesh_2_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_2_15_io_in_id_0 = r_754_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_15_io_in_id_1 = r_754_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_2_15_io_in_last_0 = r_1010_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_15_io_in_last_1 = r_1010_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_2_15_io_in_valid_0 = r_498_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_2_15_io_in_valid_1 = r_498_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_0_clock = clock;
  assign mesh_3_0_io_in_a_0 = r_48_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_0_io_in_a_1 = r_48_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_0_io_in_b_0 = pipe_b_3_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_b_1 = pipe_b_3_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_d_0 = pipe_b_259_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_d_1 = pipe_b_259_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_control_0_dataflow = mesh_3_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_control_0_propagate = mesh_3_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_control_0_shift = mesh_3_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_control_1_dataflow = mesh_3_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_control_1_propagate = mesh_3_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_control_1_shift = mesh_3_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_0_io_in_id_0 = r_515_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_0_io_in_id_1 = r_515_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_0_io_in_last_0 = r_771_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_0_io_in_last_1 = r_771_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_0_io_in_valid_0 = r_259_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_0_io_in_valid_1 = r_259_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_1_clock = clock;
  assign mesh_3_1_io_in_a_0 = r_49_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_1_io_in_a_1 = r_49_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_1_io_in_b_0 = pipe_b_19_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_b_1 = pipe_b_19_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_d_0 = pipe_b_275_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_d_1 = pipe_b_275_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_control_0_dataflow = mesh_3_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_control_0_propagate = mesh_3_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_control_0_shift = mesh_3_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_control_1_dataflow = mesh_3_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_control_1_propagate = mesh_3_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_control_1_shift = mesh_3_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_1_io_in_id_0 = r_531_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_1_io_in_id_1 = r_531_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_1_io_in_last_0 = r_787_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_1_io_in_last_1 = r_787_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_1_io_in_valid_0 = r_275_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_1_io_in_valid_1 = r_275_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_2_clock = clock;
  assign mesh_3_2_io_in_a_0 = r_50_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_2_io_in_a_1 = r_50_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_2_io_in_b_0 = pipe_b_35_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_b_1 = pipe_b_35_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_d_0 = pipe_b_291_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_d_1 = pipe_b_291_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_control_0_dataflow = mesh_3_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_control_0_propagate = mesh_3_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_control_0_shift = mesh_3_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_control_1_dataflow = mesh_3_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_control_1_propagate = mesh_3_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_control_1_shift = mesh_3_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_2_io_in_id_0 = r_547_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_2_io_in_id_1 = r_547_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_2_io_in_last_0 = r_803_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_2_io_in_last_1 = r_803_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_2_io_in_valid_0 = r_291_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_2_io_in_valid_1 = r_291_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_3_clock = clock;
  assign mesh_3_3_io_in_a_0 = r_51_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_3_io_in_a_1 = r_51_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_3_io_in_b_0 = pipe_b_51_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_b_1 = pipe_b_51_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_d_0 = pipe_b_307_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_d_1 = pipe_b_307_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_control_0_dataflow = mesh_3_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_control_0_propagate = mesh_3_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_control_0_shift = mesh_3_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_control_1_dataflow = mesh_3_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_control_1_propagate = mesh_3_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_control_1_shift = mesh_3_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_3_io_in_id_0 = r_563_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_3_io_in_id_1 = r_563_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_3_io_in_last_0 = r_819_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_3_io_in_last_1 = r_819_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_3_io_in_valid_0 = r_307_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_3_io_in_valid_1 = r_307_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_4_clock = clock;
  assign mesh_3_4_io_in_a_0 = r_52_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_4_io_in_a_1 = r_52_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_4_io_in_b_0 = pipe_b_67_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_b_1 = pipe_b_67_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_d_0 = pipe_b_323_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_d_1 = pipe_b_323_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_control_0_dataflow = mesh_3_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_control_0_propagate = mesh_3_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_control_0_shift = mesh_3_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_control_1_dataflow = mesh_3_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_control_1_propagate = mesh_3_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_control_1_shift = mesh_3_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_4_io_in_id_0 = r_579_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_4_io_in_id_1 = r_579_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_4_io_in_last_0 = r_835_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_4_io_in_last_1 = r_835_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_4_io_in_valid_0 = r_323_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_4_io_in_valid_1 = r_323_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_5_clock = clock;
  assign mesh_3_5_io_in_a_0 = r_53_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_5_io_in_a_1 = r_53_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_5_io_in_b_0 = pipe_b_83_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_b_1 = pipe_b_83_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_d_0 = pipe_b_339_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_d_1 = pipe_b_339_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_control_0_dataflow = mesh_3_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_control_0_propagate = mesh_3_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_control_0_shift = mesh_3_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_control_1_dataflow = mesh_3_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_control_1_propagate = mesh_3_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_control_1_shift = mesh_3_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_5_io_in_id_0 = r_595_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_5_io_in_id_1 = r_595_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_5_io_in_last_0 = r_851_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_5_io_in_last_1 = r_851_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_5_io_in_valid_0 = r_339_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_5_io_in_valid_1 = r_339_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_6_clock = clock;
  assign mesh_3_6_io_in_a_0 = r_54_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_6_io_in_a_1 = r_54_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_6_io_in_b_0 = pipe_b_99_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_b_1 = pipe_b_99_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_d_0 = pipe_b_355_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_d_1 = pipe_b_355_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_control_0_dataflow = mesh_3_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_control_0_propagate = mesh_3_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_control_0_shift = mesh_3_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_control_1_dataflow = mesh_3_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_control_1_propagate = mesh_3_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_control_1_shift = mesh_3_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_6_io_in_id_0 = r_611_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_6_io_in_id_1 = r_611_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_6_io_in_last_0 = r_867_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_6_io_in_last_1 = r_867_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_6_io_in_valid_0 = r_355_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_6_io_in_valid_1 = r_355_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_7_clock = clock;
  assign mesh_3_7_io_in_a_0 = r_55_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_7_io_in_a_1 = r_55_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_7_io_in_b_0 = pipe_b_115_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_b_1 = pipe_b_115_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_d_0 = pipe_b_371_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_d_1 = pipe_b_371_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_control_0_dataflow = mesh_3_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_control_0_propagate = mesh_3_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_control_0_shift = mesh_3_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_control_1_dataflow = mesh_3_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_control_1_propagate = mesh_3_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_control_1_shift = mesh_3_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_7_io_in_id_0 = r_627_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_7_io_in_id_1 = r_627_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_7_io_in_last_0 = r_883_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_7_io_in_last_1 = r_883_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_7_io_in_valid_0 = r_371_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_7_io_in_valid_1 = r_371_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_8_clock = clock;
  assign mesh_3_8_io_in_a_0 = r_56_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_8_io_in_a_1 = r_56_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_8_io_in_b_0 = pipe_b_131_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_b_1 = pipe_b_131_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_d_0 = pipe_b_387_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_d_1 = pipe_b_387_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_control_0_dataflow = mesh_3_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_control_0_propagate = mesh_3_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_control_0_shift = mesh_3_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_control_1_dataflow = mesh_3_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_control_1_propagate = mesh_3_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_control_1_shift = mesh_3_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_8_io_in_id_0 = r_643_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_8_io_in_id_1 = r_643_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_8_io_in_last_0 = r_899_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_8_io_in_last_1 = r_899_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_8_io_in_valid_0 = r_387_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_8_io_in_valid_1 = r_387_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_9_clock = clock;
  assign mesh_3_9_io_in_a_0 = r_57_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_9_io_in_a_1 = r_57_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_9_io_in_b_0 = pipe_b_147_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_b_1 = pipe_b_147_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_d_0 = pipe_b_403_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_d_1 = pipe_b_403_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_control_0_dataflow = mesh_3_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_control_0_propagate = mesh_3_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_control_0_shift = mesh_3_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_control_1_dataflow = mesh_3_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_control_1_propagate = mesh_3_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_control_1_shift = mesh_3_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_9_io_in_id_0 = r_659_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_9_io_in_id_1 = r_659_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_9_io_in_last_0 = r_915_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_9_io_in_last_1 = r_915_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_9_io_in_valid_0 = r_403_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_9_io_in_valid_1 = r_403_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_10_clock = clock;
  assign mesh_3_10_io_in_a_0 = r_58_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_10_io_in_a_1 = r_58_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_10_io_in_b_0 = pipe_b_163_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_b_1 = pipe_b_163_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_d_0 = pipe_b_419_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_d_1 = pipe_b_419_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_control_0_dataflow = mesh_3_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_control_0_propagate = mesh_3_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_control_0_shift = mesh_3_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_control_1_dataflow = mesh_3_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_control_1_propagate = mesh_3_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_control_1_shift = mesh_3_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_10_io_in_id_0 = r_675_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_10_io_in_id_1 = r_675_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_10_io_in_last_0 = r_931_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_10_io_in_last_1 = r_931_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_10_io_in_valid_0 = r_419_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_10_io_in_valid_1 = r_419_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_11_clock = clock;
  assign mesh_3_11_io_in_a_0 = r_59_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_11_io_in_a_1 = r_59_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_11_io_in_b_0 = pipe_b_179_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_b_1 = pipe_b_179_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_d_0 = pipe_b_435_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_d_1 = pipe_b_435_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_control_0_dataflow = mesh_3_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_control_0_propagate = mesh_3_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_control_0_shift = mesh_3_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_control_1_dataflow = mesh_3_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_control_1_propagate = mesh_3_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_control_1_shift = mesh_3_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_11_io_in_id_0 = r_691_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_11_io_in_id_1 = r_691_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_11_io_in_last_0 = r_947_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_11_io_in_last_1 = r_947_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_11_io_in_valid_0 = r_435_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_11_io_in_valid_1 = r_435_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_12_clock = clock;
  assign mesh_3_12_io_in_a_0 = r_60_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_12_io_in_a_1 = r_60_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_12_io_in_b_0 = pipe_b_195_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_b_1 = pipe_b_195_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_d_0 = pipe_b_451_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_d_1 = pipe_b_451_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_control_0_dataflow = mesh_3_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_control_0_propagate = mesh_3_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_control_0_shift = mesh_3_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_control_1_dataflow = mesh_3_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_control_1_propagate = mesh_3_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_control_1_shift = mesh_3_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_12_io_in_id_0 = r_707_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_12_io_in_id_1 = r_707_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_12_io_in_last_0 = r_963_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_12_io_in_last_1 = r_963_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_12_io_in_valid_0 = r_451_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_12_io_in_valid_1 = r_451_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_13_clock = clock;
  assign mesh_3_13_io_in_a_0 = r_61_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_13_io_in_a_1 = r_61_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_13_io_in_b_0 = pipe_b_211_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_b_1 = pipe_b_211_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_d_0 = pipe_b_467_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_d_1 = pipe_b_467_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_control_0_dataflow = mesh_3_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_control_0_propagate = mesh_3_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_control_0_shift = mesh_3_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_control_1_dataflow = mesh_3_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_control_1_propagate = mesh_3_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_control_1_shift = mesh_3_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_13_io_in_id_0 = r_723_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_13_io_in_id_1 = r_723_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_13_io_in_last_0 = r_979_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_13_io_in_last_1 = r_979_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_13_io_in_valid_0 = r_467_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_13_io_in_valid_1 = r_467_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_14_clock = clock;
  assign mesh_3_14_io_in_a_0 = r_62_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_14_io_in_a_1 = r_62_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_14_io_in_b_0 = pipe_b_227_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_b_1 = pipe_b_227_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_d_0 = pipe_b_483_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_d_1 = pipe_b_483_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_control_0_dataflow = mesh_3_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_control_0_propagate = mesh_3_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_control_0_shift = mesh_3_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_control_1_dataflow = mesh_3_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_control_1_propagate = mesh_3_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_control_1_shift = mesh_3_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_14_io_in_id_0 = r_739_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_14_io_in_id_1 = r_739_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_14_io_in_last_0 = r_995_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_14_io_in_last_1 = r_995_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_14_io_in_valid_0 = r_483_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_14_io_in_valid_1 = r_483_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_15_clock = clock;
  assign mesh_3_15_io_in_a_0 = r_63_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_15_io_in_a_1 = r_63_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_3_15_io_in_b_0 = pipe_b_243_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_b_1 = pipe_b_243_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_d_0 = pipe_b_499_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_d_1 = pipe_b_499_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_control_0_dataflow = mesh_3_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_control_0_propagate = mesh_3_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_control_0_shift = mesh_3_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_control_1_dataflow = mesh_3_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_control_1_propagate = mesh_3_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_control_1_shift = mesh_3_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_3_15_io_in_id_0 = r_755_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_15_io_in_id_1 = r_755_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_3_15_io_in_last_0 = r_1011_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_15_io_in_last_1 = r_1011_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_3_15_io_in_valid_0 = r_499_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_3_15_io_in_valid_1 = r_499_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_0_clock = clock;
  assign mesh_4_0_io_in_a_0 = r_64_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_0_io_in_a_1 = r_64_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_0_io_in_b_0 = pipe_b_4_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_b_1 = pipe_b_4_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_d_0 = pipe_b_260_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_d_1 = pipe_b_260_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_control_0_dataflow = mesh_4_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_control_0_propagate = mesh_4_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_control_0_shift = mesh_4_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_control_1_dataflow = mesh_4_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_control_1_propagate = mesh_4_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_control_1_shift = mesh_4_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_0_io_in_id_0 = r_516_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_0_io_in_id_1 = r_516_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_0_io_in_last_0 = r_772_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_0_io_in_last_1 = r_772_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_0_io_in_valid_0 = r_260_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_0_io_in_valid_1 = r_260_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_1_clock = clock;
  assign mesh_4_1_io_in_a_0 = r_65_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_1_io_in_a_1 = r_65_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_1_io_in_b_0 = pipe_b_20_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_b_1 = pipe_b_20_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_d_0 = pipe_b_276_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_d_1 = pipe_b_276_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_control_0_dataflow = mesh_4_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_control_0_propagate = mesh_4_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_control_0_shift = mesh_4_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_control_1_dataflow = mesh_4_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_control_1_propagate = mesh_4_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_control_1_shift = mesh_4_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_1_io_in_id_0 = r_532_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_1_io_in_id_1 = r_532_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_1_io_in_last_0 = r_788_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_1_io_in_last_1 = r_788_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_1_io_in_valid_0 = r_276_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_1_io_in_valid_1 = r_276_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_2_clock = clock;
  assign mesh_4_2_io_in_a_0 = r_66_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_2_io_in_a_1 = r_66_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_2_io_in_b_0 = pipe_b_36_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_b_1 = pipe_b_36_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_d_0 = pipe_b_292_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_d_1 = pipe_b_292_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_control_0_dataflow = mesh_4_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_control_0_propagate = mesh_4_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_control_0_shift = mesh_4_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_control_1_dataflow = mesh_4_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_control_1_propagate = mesh_4_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_control_1_shift = mesh_4_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_2_io_in_id_0 = r_548_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_2_io_in_id_1 = r_548_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_2_io_in_last_0 = r_804_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_2_io_in_last_1 = r_804_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_2_io_in_valid_0 = r_292_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_2_io_in_valid_1 = r_292_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_3_clock = clock;
  assign mesh_4_3_io_in_a_0 = r_67_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_3_io_in_a_1 = r_67_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_3_io_in_b_0 = pipe_b_52_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_b_1 = pipe_b_52_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_d_0 = pipe_b_308_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_d_1 = pipe_b_308_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_control_0_dataflow = mesh_4_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_control_0_propagate = mesh_4_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_control_0_shift = mesh_4_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_control_1_dataflow = mesh_4_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_control_1_propagate = mesh_4_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_control_1_shift = mesh_4_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_3_io_in_id_0 = r_564_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_3_io_in_id_1 = r_564_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_3_io_in_last_0 = r_820_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_3_io_in_last_1 = r_820_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_3_io_in_valid_0 = r_308_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_3_io_in_valid_1 = r_308_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_4_clock = clock;
  assign mesh_4_4_io_in_a_0 = r_68_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_4_io_in_a_1 = r_68_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_4_io_in_b_0 = pipe_b_68_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_b_1 = pipe_b_68_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_d_0 = pipe_b_324_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_d_1 = pipe_b_324_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_control_0_dataflow = mesh_4_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_control_0_propagate = mesh_4_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_control_0_shift = mesh_4_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_control_1_dataflow = mesh_4_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_control_1_propagate = mesh_4_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_control_1_shift = mesh_4_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_4_io_in_id_0 = r_580_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_4_io_in_id_1 = r_580_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_4_io_in_last_0 = r_836_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_4_io_in_last_1 = r_836_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_4_io_in_valid_0 = r_324_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_4_io_in_valid_1 = r_324_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_5_clock = clock;
  assign mesh_4_5_io_in_a_0 = r_69_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_5_io_in_a_1 = r_69_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_5_io_in_b_0 = pipe_b_84_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_b_1 = pipe_b_84_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_d_0 = pipe_b_340_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_d_1 = pipe_b_340_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_control_0_dataflow = mesh_4_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_control_0_propagate = mesh_4_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_control_0_shift = mesh_4_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_control_1_dataflow = mesh_4_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_control_1_propagate = mesh_4_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_control_1_shift = mesh_4_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_5_io_in_id_0 = r_596_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_5_io_in_id_1 = r_596_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_5_io_in_last_0 = r_852_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_5_io_in_last_1 = r_852_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_5_io_in_valid_0 = r_340_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_5_io_in_valid_1 = r_340_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_6_clock = clock;
  assign mesh_4_6_io_in_a_0 = r_70_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_6_io_in_a_1 = r_70_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_6_io_in_b_0 = pipe_b_100_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_b_1 = pipe_b_100_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_d_0 = pipe_b_356_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_d_1 = pipe_b_356_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_control_0_dataflow = mesh_4_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_control_0_propagate = mesh_4_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_control_0_shift = mesh_4_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_control_1_dataflow = mesh_4_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_control_1_propagate = mesh_4_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_control_1_shift = mesh_4_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_6_io_in_id_0 = r_612_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_6_io_in_id_1 = r_612_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_6_io_in_last_0 = r_868_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_6_io_in_last_1 = r_868_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_6_io_in_valid_0 = r_356_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_6_io_in_valid_1 = r_356_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_7_clock = clock;
  assign mesh_4_7_io_in_a_0 = r_71_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_7_io_in_a_1 = r_71_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_7_io_in_b_0 = pipe_b_116_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_b_1 = pipe_b_116_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_d_0 = pipe_b_372_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_d_1 = pipe_b_372_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_control_0_dataflow = mesh_4_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_control_0_propagate = mesh_4_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_control_0_shift = mesh_4_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_control_1_dataflow = mesh_4_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_control_1_propagate = mesh_4_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_control_1_shift = mesh_4_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_7_io_in_id_0 = r_628_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_7_io_in_id_1 = r_628_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_7_io_in_last_0 = r_884_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_7_io_in_last_1 = r_884_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_7_io_in_valid_0 = r_372_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_7_io_in_valid_1 = r_372_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_8_clock = clock;
  assign mesh_4_8_io_in_a_0 = r_72_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_8_io_in_a_1 = r_72_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_8_io_in_b_0 = pipe_b_132_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_b_1 = pipe_b_132_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_d_0 = pipe_b_388_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_d_1 = pipe_b_388_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_control_0_dataflow = mesh_4_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_control_0_propagate = mesh_4_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_control_0_shift = mesh_4_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_control_1_dataflow = mesh_4_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_control_1_propagate = mesh_4_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_control_1_shift = mesh_4_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_8_io_in_id_0 = r_644_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_8_io_in_id_1 = r_644_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_8_io_in_last_0 = r_900_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_8_io_in_last_1 = r_900_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_8_io_in_valid_0 = r_388_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_8_io_in_valid_1 = r_388_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_9_clock = clock;
  assign mesh_4_9_io_in_a_0 = r_73_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_9_io_in_a_1 = r_73_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_9_io_in_b_0 = pipe_b_148_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_b_1 = pipe_b_148_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_d_0 = pipe_b_404_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_d_1 = pipe_b_404_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_control_0_dataflow = mesh_4_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_control_0_propagate = mesh_4_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_control_0_shift = mesh_4_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_control_1_dataflow = mesh_4_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_control_1_propagate = mesh_4_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_control_1_shift = mesh_4_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_9_io_in_id_0 = r_660_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_9_io_in_id_1 = r_660_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_9_io_in_last_0 = r_916_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_9_io_in_last_1 = r_916_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_9_io_in_valid_0 = r_404_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_9_io_in_valid_1 = r_404_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_10_clock = clock;
  assign mesh_4_10_io_in_a_0 = r_74_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_10_io_in_a_1 = r_74_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_10_io_in_b_0 = pipe_b_164_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_b_1 = pipe_b_164_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_d_0 = pipe_b_420_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_d_1 = pipe_b_420_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_control_0_dataflow = mesh_4_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_control_0_propagate = mesh_4_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_control_0_shift = mesh_4_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_control_1_dataflow = mesh_4_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_control_1_propagate = mesh_4_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_control_1_shift = mesh_4_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_10_io_in_id_0 = r_676_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_10_io_in_id_1 = r_676_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_10_io_in_last_0 = r_932_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_10_io_in_last_1 = r_932_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_10_io_in_valid_0 = r_420_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_10_io_in_valid_1 = r_420_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_11_clock = clock;
  assign mesh_4_11_io_in_a_0 = r_75_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_11_io_in_a_1 = r_75_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_11_io_in_b_0 = pipe_b_180_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_b_1 = pipe_b_180_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_d_0 = pipe_b_436_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_d_1 = pipe_b_436_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_control_0_dataflow = mesh_4_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_control_0_propagate = mesh_4_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_control_0_shift = mesh_4_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_control_1_dataflow = mesh_4_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_control_1_propagate = mesh_4_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_control_1_shift = mesh_4_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_11_io_in_id_0 = r_692_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_11_io_in_id_1 = r_692_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_11_io_in_last_0 = r_948_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_11_io_in_last_1 = r_948_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_11_io_in_valid_0 = r_436_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_11_io_in_valid_1 = r_436_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_12_clock = clock;
  assign mesh_4_12_io_in_a_0 = r_76_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_12_io_in_a_1 = r_76_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_12_io_in_b_0 = pipe_b_196_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_b_1 = pipe_b_196_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_d_0 = pipe_b_452_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_d_1 = pipe_b_452_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_control_0_dataflow = mesh_4_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_control_0_propagate = mesh_4_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_control_0_shift = mesh_4_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_control_1_dataflow = mesh_4_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_control_1_propagate = mesh_4_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_control_1_shift = mesh_4_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_12_io_in_id_0 = r_708_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_12_io_in_id_1 = r_708_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_12_io_in_last_0 = r_964_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_12_io_in_last_1 = r_964_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_12_io_in_valid_0 = r_452_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_12_io_in_valid_1 = r_452_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_13_clock = clock;
  assign mesh_4_13_io_in_a_0 = r_77_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_13_io_in_a_1 = r_77_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_13_io_in_b_0 = pipe_b_212_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_b_1 = pipe_b_212_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_d_0 = pipe_b_468_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_d_1 = pipe_b_468_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_control_0_dataflow = mesh_4_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_control_0_propagate = mesh_4_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_control_0_shift = mesh_4_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_control_1_dataflow = mesh_4_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_control_1_propagate = mesh_4_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_control_1_shift = mesh_4_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_13_io_in_id_0 = r_724_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_13_io_in_id_1 = r_724_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_13_io_in_last_0 = r_980_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_13_io_in_last_1 = r_980_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_13_io_in_valid_0 = r_468_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_13_io_in_valid_1 = r_468_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_14_clock = clock;
  assign mesh_4_14_io_in_a_0 = r_78_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_14_io_in_a_1 = r_78_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_14_io_in_b_0 = pipe_b_228_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_b_1 = pipe_b_228_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_d_0 = pipe_b_484_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_d_1 = pipe_b_484_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_control_0_dataflow = mesh_4_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_control_0_propagate = mesh_4_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_control_0_shift = mesh_4_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_control_1_dataflow = mesh_4_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_control_1_propagate = mesh_4_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_control_1_shift = mesh_4_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_14_io_in_id_0 = r_740_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_14_io_in_id_1 = r_740_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_14_io_in_last_0 = r_996_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_14_io_in_last_1 = r_996_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_14_io_in_valid_0 = r_484_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_14_io_in_valid_1 = r_484_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_15_clock = clock;
  assign mesh_4_15_io_in_a_0 = r_79_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_15_io_in_a_1 = r_79_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_4_15_io_in_b_0 = pipe_b_244_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_b_1 = pipe_b_244_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_d_0 = pipe_b_500_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_d_1 = pipe_b_500_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_control_0_dataflow = mesh_4_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_control_0_propagate = mesh_4_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_control_0_shift = mesh_4_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_control_1_dataflow = mesh_4_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_control_1_propagate = mesh_4_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_control_1_shift = mesh_4_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_4_15_io_in_id_0 = r_756_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_15_io_in_id_1 = r_756_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_4_15_io_in_last_0 = r_1012_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_15_io_in_last_1 = r_1012_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_4_15_io_in_valid_0 = r_500_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_4_15_io_in_valid_1 = r_500_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_0_clock = clock;
  assign mesh_5_0_io_in_a_0 = r_80_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_0_io_in_a_1 = r_80_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_0_io_in_b_0 = pipe_b_5_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_b_1 = pipe_b_5_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_d_0 = pipe_b_261_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_d_1 = pipe_b_261_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_control_0_dataflow = mesh_5_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_control_0_propagate = mesh_5_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_control_0_shift = mesh_5_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_control_1_dataflow = mesh_5_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_control_1_propagate = mesh_5_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_control_1_shift = mesh_5_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_0_io_in_id_0 = r_517_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_0_io_in_id_1 = r_517_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_0_io_in_last_0 = r_773_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_0_io_in_last_1 = r_773_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_0_io_in_valid_0 = r_261_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_0_io_in_valid_1 = r_261_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_1_clock = clock;
  assign mesh_5_1_io_in_a_0 = r_81_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_1_io_in_a_1 = r_81_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_1_io_in_b_0 = pipe_b_21_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_b_1 = pipe_b_21_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_d_0 = pipe_b_277_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_d_1 = pipe_b_277_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_control_0_dataflow = mesh_5_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_control_0_propagate = mesh_5_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_control_0_shift = mesh_5_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_control_1_dataflow = mesh_5_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_control_1_propagate = mesh_5_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_control_1_shift = mesh_5_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_1_io_in_id_0 = r_533_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_1_io_in_id_1 = r_533_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_1_io_in_last_0 = r_789_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_1_io_in_last_1 = r_789_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_1_io_in_valid_0 = r_277_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_1_io_in_valid_1 = r_277_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_2_clock = clock;
  assign mesh_5_2_io_in_a_0 = r_82_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_2_io_in_a_1 = r_82_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_2_io_in_b_0 = pipe_b_37_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_b_1 = pipe_b_37_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_d_0 = pipe_b_293_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_d_1 = pipe_b_293_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_control_0_dataflow = mesh_5_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_control_0_propagate = mesh_5_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_control_0_shift = mesh_5_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_control_1_dataflow = mesh_5_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_control_1_propagate = mesh_5_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_control_1_shift = mesh_5_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_2_io_in_id_0 = r_549_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_2_io_in_id_1 = r_549_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_2_io_in_last_0 = r_805_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_2_io_in_last_1 = r_805_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_2_io_in_valid_0 = r_293_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_2_io_in_valid_1 = r_293_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_3_clock = clock;
  assign mesh_5_3_io_in_a_0 = r_83_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_3_io_in_a_1 = r_83_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_3_io_in_b_0 = pipe_b_53_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_b_1 = pipe_b_53_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_d_0 = pipe_b_309_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_d_1 = pipe_b_309_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_control_0_dataflow = mesh_5_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_control_0_propagate = mesh_5_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_control_0_shift = mesh_5_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_control_1_dataflow = mesh_5_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_control_1_propagate = mesh_5_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_control_1_shift = mesh_5_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_3_io_in_id_0 = r_565_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_3_io_in_id_1 = r_565_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_3_io_in_last_0 = r_821_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_3_io_in_last_1 = r_821_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_3_io_in_valid_0 = r_309_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_3_io_in_valid_1 = r_309_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_4_clock = clock;
  assign mesh_5_4_io_in_a_0 = r_84_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_4_io_in_a_1 = r_84_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_4_io_in_b_0 = pipe_b_69_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_b_1 = pipe_b_69_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_d_0 = pipe_b_325_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_d_1 = pipe_b_325_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_control_0_dataflow = mesh_5_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_control_0_propagate = mesh_5_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_control_0_shift = mesh_5_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_control_1_dataflow = mesh_5_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_control_1_propagate = mesh_5_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_control_1_shift = mesh_5_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_4_io_in_id_0 = r_581_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_4_io_in_id_1 = r_581_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_4_io_in_last_0 = r_837_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_4_io_in_last_1 = r_837_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_4_io_in_valid_0 = r_325_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_4_io_in_valid_1 = r_325_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_5_clock = clock;
  assign mesh_5_5_io_in_a_0 = r_85_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_5_io_in_a_1 = r_85_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_5_io_in_b_0 = pipe_b_85_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_b_1 = pipe_b_85_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_d_0 = pipe_b_341_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_d_1 = pipe_b_341_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_control_0_dataflow = mesh_5_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_control_0_propagate = mesh_5_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_control_0_shift = mesh_5_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_control_1_dataflow = mesh_5_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_control_1_propagate = mesh_5_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_control_1_shift = mesh_5_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_5_io_in_id_0 = r_597_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_5_io_in_id_1 = r_597_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_5_io_in_last_0 = r_853_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_5_io_in_last_1 = r_853_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_5_io_in_valid_0 = r_341_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_5_io_in_valid_1 = r_341_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_6_clock = clock;
  assign mesh_5_6_io_in_a_0 = r_86_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_6_io_in_a_1 = r_86_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_6_io_in_b_0 = pipe_b_101_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_b_1 = pipe_b_101_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_d_0 = pipe_b_357_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_d_1 = pipe_b_357_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_control_0_dataflow = mesh_5_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_control_0_propagate = mesh_5_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_control_0_shift = mesh_5_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_control_1_dataflow = mesh_5_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_control_1_propagate = mesh_5_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_control_1_shift = mesh_5_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_6_io_in_id_0 = r_613_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_6_io_in_id_1 = r_613_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_6_io_in_last_0 = r_869_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_6_io_in_last_1 = r_869_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_6_io_in_valid_0 = r_357_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_6_io_in_valid_1 = r_357_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_7_clock = clock;
  assign mesh_5_7_io_in_a_0 = r_87_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_7_io_in_a_1 = r_87_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_7_io_in_b_0 = pipe_b_117_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_b_1 = pipe_b_117_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_d_0 = pipe_b_373_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_d_1 = pipe_b_373_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_control_0_dataflow = mesh_5_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_control_0_propagate = mesh_5_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_control_0_shift = mesh_5_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_control_1_dataflow = mesh_5_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_control_1_propagate = mesh_5_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_control_1_shift = mesh_5_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_7_io_in_id_0 = r_629_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_7_io_in_id_1 = r_629_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_7_io_in_last_0 = r_885_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_7_io_in_last_1 = r_885_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_7_io_in_valid_0 = r_373_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_7_io_in_valid_1 = r_373_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_8_clock = clock;
  assign mesh_5_8_io_in_a_0 = r_88_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_8_io_in_a_1 = r_88_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_8_io_in_b_0 = pipe_b_133_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_b_1 = pipe_b_133_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_d_0 = pipe_b_389_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_d_1 = pipe_b_389_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_control_0_dataflow = mesh_5_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_control_0_propagate = mesh_5_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_control_0_shift = mesh_5_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_control_1_dataflow = mesh_5_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_control_1_propagate = mesh_5_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_control_1_shift = mesh_5_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_8_io_in_id_0 = r_645_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_8_io_in_id_1 = r_645_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_8_io_in_last_0 = r_901_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_8_io_in_last_1 = r_901_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_8_io_in_valid_0 = r_389_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_8_io_in_valid_1 = r_389_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_9_clock = clock;
  assign mesh_5_9_io_in_a_0 = r_89_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_9_io_in_a_1 = r_89_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_9_io_in_b_0 = pipe_b_149_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_b_1 = pipe_b_149_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_d_0 = pipe_b_405_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_d_1 = pipe_b_405_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_control_0_dataflow = mesh_5_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_control_0_propagate = mesh_5_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_control_0_shift = mesh_5_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_control_1_dataflow = mesh_5_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_control_1_propagate = mesh_5_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_control_1_shift = mesh_5_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_9_io_in_id_0 = r_661_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_9_io_in_id_1 = r_661_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_9_io_in_last_0 = r_917_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_9_io_in_last_1 = r_917_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_9_io_in_valid_0 = r_405_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_9_io_in_valid_1 = r_405_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_10_clock = clock;
  assign mesh_5_10_io_in_a_0 = r_90_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_10_io_in_a_1 = r_90_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_10_io_in_b_0 = pipe_b_165_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_b_1 = pipe_b_165_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_d_0 = pipe_b_421_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_d_1 = pipe_b_421_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_control_0_dataflow = mesh_5_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_control_0_propagate = mesh_5_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_control_0_shift = mesh_5_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_control_1_dataflow = mesh_5_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_control_1_propagate = mesh_5_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_control_1_shift = mesh_5_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_10_io_in_id_0 = r_677_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_10_io_in_id_1 = r_677_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_10_io_in_last_0 = r_933_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_10_io_in_last_1 = r_933_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_10_io_in_valid_0 = r_421_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_10_io_in_valid_1 = r_421_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_11_clock = clock;
  assign mesh_5_11_io_in_a_0 = r_91_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_11_io_in_a_1 = r_91_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_11_io_in_b_0 = pipe_b_181_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_b_1 = pipe_b_181_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_d_0 = pipe_b_437_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_d_1 = pipe_b_437_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_control_0_dataflow = mesh_5_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_control_0_propagate = mesh_5_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_control_0_shift = mesh_5_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_control_1_dataflow = mesh_5_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_control_1_propagate = mesh_5_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_control_1_shift = mesh_5_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_11_io_in_id_0 = r_693_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_11_io_in_id_1 = r_693_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_11_io_in_last_0 = r_949_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_11_io_in_last_1 = r_949_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_11_io_in_valid_0 = r_437_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_11_io_in_valid_1 = r_437_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_12_clock = clock;
  assign mesh_5_12_io_in_a_0 = r_92_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_12_io_in_a_1 = r_92_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_12_io_in_b_0 = pipe_b_197_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_b_1 = pipe_b_197_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_d_0 = pipe_b_453_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_d_1 = pipe_b_453_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_control_0_dataflow = mesh_5_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_control_0_propagate = mesh_5_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_control_0_shift = mesh_5_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_control_1_dataflow = mesh_5_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_control_1_propagate = mesh_5_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_control_1_shift = mesh_5_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_12_io_in_id_0 = r_709_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_12_io_in_id_1 = r_709_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_12_io_in_last_0 = r_965_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_12_io_in_last_1 = r_965_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_12_io_in_valid_0 = r_453_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_12_io_in_valid_1 = r_453_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_13_clock = clock;
  assign mesh_5_13_io_in_a_0 = r_93_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_13_io_in_a_1 = r_93_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_13_io_in_b_0 = pipe_b_213_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_b_1 = pipe_b_213_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_d_0 = pipe_b_469_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_d_1 = pipe_b_469_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_control_0_dataflow = mesh_5_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_control_0_propagate = mesh_5_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_control_0_shift = mesh_5_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_control_1_dataflow = mesh_5_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_control_1_propagate = mesh_5_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_control_1_shift = mesh_5_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_13_io_in_id_0 = r_725_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_13_io_in_id_1 = r_725_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_13_io_in_last_0 = r_981_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_13_io_in_last_1 = r_981_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_13_io_in_valid_0 = r_469_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_13_io_in_valid_1 = r_469_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_14_clock = clock;
  assign mesh_5_14_io_in_a_0 = r_94_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_14_io_in_a_1 = r_94_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_14_io_in_b_0 = pipe_b_229_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_b_1 = pipe_b_229_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_d_0 = pipe_b_485_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_d_1 = pipe_b_485_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_control_0_dataflow = mesh_5_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_control_0_propagate = mesh_5_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_control_0_shift = mesh_5_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_control_1_dataflow = mesh_5_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_control_1_propagate = mesh_5_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_control_1_shift = mesh_5_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_14_io_in_id_0 = r_741_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_14_io_in_id_1 = r_741_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_14_io_in_last_0 = r_997_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_14_io_in_last_1 = r_997_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_14_io_in_valid_0 = r_485_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_14_io_in_valid_1 = r_485_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_15_clock = clock;
  assign mesh_5_15_io_in_a_0 = r_95_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_15_io_in_a_1 = r_95_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_5_15_io_in_b_0 = pipe_b_245_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_b_1 = pipe_b_245_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_d_0 = pipe_b_501_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_d_1 = pipe_b_501_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_control_0_dataflow = mesh_5_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_control_0_propagate = mesh_5_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_control_0_shift = mesh_5_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_control_1_dataflow = mesh_5_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_control_1_propagate = mesh_5_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_control_1_shift = mesh_5_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_5_15_io_in_id_0 = r_757_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_15_io_in_id_1 = r_757_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_5_15_io_in_last_0 = r_1013_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_15_io_in_last_1 = r_1013_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_5_15_io_in_valid_0 = r_501_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_5_15_io_in_valid_1 = r_501_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_0_clock = clock;
  assign mesh_6_0_io_in_a_0 = r_96_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_0_io_in_a_1 = r_96_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_0_io_in_b_0 = pipe_b_6_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_b_1 = pipe_b_6_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_d_0 = pipe_b_262_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_d_1 = pipe_b_262_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_control_0_dataflow = mesh_6_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_control_0_propagate = mesh_6_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_control_0_shift = mesh_6_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_control_1_dataflow = mesh_6_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_control_1_propagate = mesh_6_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_control_1_shift = mesh_6_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_0_io_in_id_0 = r_518_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_0_io_in_id_1 = r_518_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_0_io_in_last_0 = r_774_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_0_io_in_last_1 = r_774_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_0_io_in_valid_0 = r_262_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_0_io_in_valid_1 = r_262_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_1_clock = clock;
  assign mesh_6_1_io_in_a_0 = r_97_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_1_io_in_a_1 = r_97_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_1_io_in_b_0 = pipe_b_22_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_b_1 = pipe_b_22_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_d_0 = pipe_b_278_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_d_1 = pipe_b_278_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_control_0_dataflow = mesh_6_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_control_0_propagate = mesh_6_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_control_0_shift = mesh_6_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_control_1_dataflow = mesh_6_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_control_1_propagate = mesh_6_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_control_1_shift = mesh_6_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_1_io_in_id_0 = r_534_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_1_io_in_id_1 = r_534_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_1_io_in_last_0 = r_790_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_1_io_in_last_1 = r_790_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_1_io_in_valid_0 = r_278_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_1_io_in_valid_1 = r_278_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_2_clock = clock;
  assign mesh_6_2_io_in_a_0 = r_98_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_2_io_in_a_1 = r_98_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_2_io_in_b_0 = pipe_b_38_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_b_1 = pipe_b_38_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_d_0 = pipe_b_294_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_d_1 = pipe_b_294_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_control_0_dataflow = mesh_6_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_control_0_propagate = mesh_6_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_control_0_shift = mesh_6_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_control_1_dataflow = mesh_6_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_control_1_propagate = mesh_6_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_control_1_shift = mesh_6_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_2_io_in_id_0 = r_550_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_2_io_in_id_1 = r_550_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_2_io_in_last_0 = r_806_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_2_io_in_last_1 = r_806_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_2_io_in_valid_0 = r_294_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_2_io_in_valid_1 = r_294_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_3_clock = clock;
  assign mesh_6_3_io_in_a_0 = r_99_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_3_io_in_a_1 = r_99_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_3_io_in_b_0 = pipe_b_54_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_b_1 = pipe_b_54_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_d_0 = pipe_b_310_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_d_1 = pipe_b_310_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_control_0_dataflow = mesh_6_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_control_0_propagate = mesh_6_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_control_0_shift = mesh_6_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_control_1_dataflow = mesh_6_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_control_1_propagate = mesh_6_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_control_1_shift = mesh_6_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_3_io_in_id_0 = r_566_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_3_io_in_id_1 = r_566_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_3_io_in_last_0 = r_822_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_3_io_in_last_1 = r_822_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_3_io_in_valid_0 = r_310_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_3_io_in_valid_1 = r_310_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_4_clock = clock;
  assign mesh_6_4_io_in_a_0 = r_100_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_4_io_in_a_1 = r_100_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_4_io_in_b_0 = pipe_b_70_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_b_1 = pipe_b_70_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_d_0 = pipe_b_326_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_d_1 = pipe_b_326_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_control_0_dataflow = mesh_6_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_control_0_propagate = mesh_6_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_control_0_shift = mesh_6_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_control_1_dataflow = mesh_6_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_control_1_propagate = mesh_6_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_control_1_shift = mesh_6_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_4_io_in_id_0 = r_582_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_4_io_in_id_1 = r_582_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_4_io_in_last_0 = r_838_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_4_io_in_last_1 = r_838_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_4_io_in_valid_0 = r_326_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_4_io_in_valid_1 = r_326_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_5_clock = clock;
  assign mesh_6_5_io_in_a_0 = r_101_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_5_io_in_a_1 = r_101_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_5_io_in_b_0 = pipe_b_86_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_b_1 = pipe_b_86_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_d_0 = pipe_b_342_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_d_1 = pipe_b_342_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_control_0_dataflow = mesh_6_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_control_0_propagate = mesh_6_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_control_0_shift = mesh_6_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_control_1_dataflow = mesh_6_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_control_1_propagate = mesh_6_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_control_1_shift = mesh_6_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_5_io_in_id_0 = r_598_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_5_io_in_id_1 = r_598_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_5_io_in_last_0 = r_854_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_5_io_in_last_1 = r_854_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_5_io_in_valid_0 = r_342_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_5_io_in_valid_1 = r_342_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_6_clock = clock;
  assign mesh_6_6_io_in_a_0 = r_102_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_6_io_in_a_1 = r_102_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_6_io_in_b_0 = pipe_b_102_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_b_1 = pipe_b_102_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_d_0 = pipe_b_358_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_d_1 = pipe_b_358_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_control_0_dataflow = mesh_6_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_control_0_propagate = mesh_6_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_control_0_shift = mesh_6_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_control_1_dataflow = mesh_6_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_control_1_propagate = mesh_6_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_control_1_shift = mesh_6_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_6_io_in_id_0 = r_614_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_6_io_in_id_1 = r_614_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_6_io_in_last_0 = r_870_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_6_io_in_last_1 = r_870_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_6_io_in_valid_0 = r_358_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_6_io_in_valid_1 = r_358_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_7_clock = clock;
  assign mesh_6_7_io_in_a_0 = r_103_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_7_io_in_a_1 = r_103_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_7_io_in_b_0 = pipe_b_118_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_b_1 = pipe_b_118_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_d_0 = pipe_b_374_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_d_1 = pipe_b_374_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_control_0_dataflow = mesh_6_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_control_0_propagate = mesh_6_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_control_0_shift = mesh_6_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_control_1_dataflow = mesh_6_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_control_1_propagate = mesh_6_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_control_1_shift = mesh_6_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_7_io_in_id_0 = r_630_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_7_io_in_id_1 = r_630_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_7_io_in_last_0 = r_886_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_7_io_in_last_1 = r_886_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_7_io_in_valid_0 = r_374_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_7_io_in_valid_1 = r_374_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_8_clock = clock;
  assign mesh_6_8_io_in_a_0 = r_104_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_8_io_in_a_1 = r_104_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_8_io_in_b_0 = pipe_b_134_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_b_1 = pipe_b_134_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_d_0 = pipe_b_390_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_d_1 = pipe_b_390_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_control_0_dataflow = mesh_6_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_control_0_propagate = mesh_6_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_control_0_shift = mesh_6_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_control_1_dataflow = mesh_6_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_control_1_propagate = mesh_6_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_control_1_shift = mesh_6_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_8_io_in_id_0 = r_646_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_8_io_in_id_1 = r_646_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_8_io_in_last_0 = r_902_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_8_io_in_last_1 = r_902_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_8_io_in_valid_0 = r_390_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_8_io_in_valid_1 = r_390_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_9_clock = clock;
  assign mesh_6_9_io_in_a_0 = r_105_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_9_io_in_a_1 = r_105_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_9_io_in_b_0 = pipe_b_150_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_b_1 = pipe_b_150_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_d_0 = pipe_b_406_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_d_1 = pipe_b_406_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_control_0_dataflow = mesh_6_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_control_0_propagate = mesh_6_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_control_0_shift = mesh_6_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_control_1_dataflow = mesh_6_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_control_1_propagate = mesh_6_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_control_1_shift = mesh_6_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_9_io_in_id_0 = r_662_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_9_io_in_id_1 = r_662_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_9_io_in_last_0 = r_918_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_9_io_in_last_1 = r_918_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_9_io_in_valid_0 = r_406_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_9_io_in_valid_1 = r_406_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_10_clock = clock;
  assign mesh_6_10_io_in_a_0 = r_106_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_10_io_in_a_1 = r_106_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_10_io_in_b_0 = pipe_b_166_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_b_1 = pipe_b_166_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_d_0 = pipe_b_422_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_d_1 = pipe_b_422_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_control_0_dataflow = mesh_6_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_control_0_propagate = mesh_6_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_control_0_shift = mesh_6_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_control_1_dataflow = mesh_6_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_control_1_propagate = mesh_6_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_control_1_shift = mesh_6_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_10_io_in_id_0 = r_678_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_10_io_in_id_1 = r_678_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_10_io_in_last_0 = r_934_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_10_io_in_last_1 = r_934_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_10_io_in_valid_0 = r_422_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_10_io_in_valid_1 = r_422_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_11_clock = clock;
  assign mesh_6_11_io_in_a_0 = r_107_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_11_io_in_a_1 = r_107_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_11_io_in_b_0 = pipe_b_182_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_b_1 = pipe_b_182_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_d_0 = pipe_b_438_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_d_1 = pipe_b_438_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_control_0_dataflow = mesh_6_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_control_0_propagate = mesh_6_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_control_0_shift = mesh_6_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_control_1_dataflow = mesh_6_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_control_1_propagate = mesh_6_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_control_1_shift = mesh_6_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_11_io_in_id_0 = r_694_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_11_io_in_id_1 = r_694_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_11_io_in_last_0 = r_950_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_11_io_in_last_1 = r_950_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_11_io_in_valid_0 = r_438_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_11_io_in_valid_1 = r_438_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_12_clock = clock;
  assign mesh_6_12_io_in_a_0 = r_108_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_12_io_in_a_1 = r_108_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_12_io_in_b_0 = pipe_b_198_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_b_1 = pipe_b_198_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_d_0 = pipe_b_454_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_d_1 = pipe_b_454_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_control_0_dataflow = mesh_6_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_control_0_propagate = mesh_6_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_control_0_shift = mesh_6_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_control_1_dataflow = mesh_6_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_control_1_propagate = mesh_6_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_control_1_shift = mesh_6_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_12_io_in_id_0 = r_710_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_12_io_in_id_1 = r_710_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_12_io_in_last_0 = r_966_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_12_io_in_last_1 = r_966_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_12_io_in_valid_0 = r_454_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_12_io_in_valid_1 = r_454_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_13_clock = clock;
  assign mesh_6_13_io_in_a_0 = r_109_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_13_io_in_a_1 = r_109_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_13_io_in_b_0 = pipe_b_214_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_b_1 = pipe_b_214_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_d_0 = pipe_b_470_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_d_1 = pipe_b_470_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_control_0_dataflow = mesh_6_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_control_0_propagate = mesh_6_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_control_0_shift = mesh_6_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_control_1_dataflow = mesh_6_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_control_1_propagate = mesh_6_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_control_1_shift = mesh_6_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_13_io_in_id_0 = r_726_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_13_io_in_id_1 = r_726_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_13_io_in_last_0 = r_982_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_13_io_in_last_1 = r_982_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_13_io_in_valid_0 = r_470_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_13_io_in_valid_1 = r_470_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_14_clock = clock;
  assign mesh_6_14_io_in_a_0 = r_110_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_14_io_in_a_1 = r_110_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_14_io_in_b_0 = pipe_b_230_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_b_1 = pipe_b_230_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_d_0 = pipe_b_486_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_d_1 = pipe_b_486_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_control_0_dataflow = mesh_6_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_control_0_propagate = mesh_6_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_control_0_shift = mesh_6_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_control_1_dataflow = mesh_6_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_control_1_propagate = mesh_6_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_control_1_shift = mesh_6_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_14_io_in_id_0 = r_742_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_14_io_in_id_1 = r_742_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_14_io_in_last_0 = r_998_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_14_io_in_last_1 = r_998_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_14_io_in_valid_0 = r_486_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_14_io_in_valid_1 = r_486_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_15_clock = clock;
  assign mesh_6_15_io_in_a_0 = r_111_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_15_io_in_a_1 = r_111_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_6_15_io_in_b_0 = pipe_b_246_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_b_1 = pipe_b_246_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_d_0 = pipe_b_502_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_d_1 = pipe_b_502_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_control_0_dataflow = mesh_6_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_control_0_propagate = mesh_6_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_control_0_shift = mesh_6_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_control_1_dataflow = mesh_6_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_control_1_propagate = mesh_6_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_control_1_shift = mesh_6_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_6_15_io_in_id_0 = r_758_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_15_io_in_id_1 = r_758_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_6_15_io_in_last_0 = r_1014_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_15_io_in_last_1 = r_1014_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_6_15_io_in_valid_0 = r_502_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_6_15_io_in_valid_1 = r_502_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_0_clock = clock;
  assign mesh_7_0_io_in_a_0 = r_112_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_0_io_in_a_1 = r_112_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_0_io_in_b_0 = pipe_b_7_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_b_1 = pipe_b_7_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_d_0 = pipe_b_263_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_d_1 = pipe_b_263_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_control_0_dataflow = mesh_7_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_control_0_propagate = mesh_7_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_control_0_shift = mesh_7_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_control_1_dataflow = mesh_7_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_control_1_propagate = mesh_7_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_control_1_shift = mesh_7_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_0_io_in_id_0 = r_519_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_0_io_in_id_1 = r_519_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_0_io_in_last_0 = r_775_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_0_io_in_last_1 = r_775_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_0_io_in_valid_0 = r_263_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_0_io_in_valid_1 = r_263_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_1_clock = clock;
  assign mesh_7_1_io_in_a_0 = r_113_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_1_io_in_a_1 = r_113_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_1_io_in_b_0 = pipe_b_23_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_b_1 = pipe_b_23_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_d_0 = pipe_b_279_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_d_1 = pipe_b_279_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_control_0_dataflow = mesh_7_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_control_0_propagate = mesh_7_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_control_0_shift = mesh_7_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_control_1_dataflow = mesh_7_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_control_1_propagate = mesh_7_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_control_1_shift = mesh_7_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_1_io_in_id_0 = r_535_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_1_io_in_id_1 = r_535_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_1_io_in_last_0 = r_791_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_1_io_in_last_1 = r_791_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_1_io_in_valid_0 = r_279_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_1_io_in_valid_1 = r_279_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_2_clock = clock;
  assign mesh_7_2_io_in_a_0 = r_114_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_2_io_in_a_1 = r_114_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_2_io_in_b_0 = pipe_b_39_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_b_1 = pipe_b_39_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_d_0 = pipe_b_295_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_d_1 = pipe_b_295_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_control_0_dataflow = mesh_7_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_control_0_propagate = mesh_7_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_control_0_shift = mesh_7_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_control_1_dataflow = mesh_7_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_control_1_propagate = mesh_7_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_control_1_shift = mesh_7_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_2_io_in_id_0 = r_551_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_2_io_in_id_1 = r_551_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_2_io_in_last_0 = r_807_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_2_io_in_last_1 = r_807_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_2_io_in_valid_0 = r_295_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_2_io_in_valid_1 = r_295_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_3_clock = clock;
  assign mesh_7_3_io_in_a_0 = r_115_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_3_io_in_a_1 = r_115_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_3_io_in_b_0 = pipe_b_55_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_b_1 = pipe_b_55_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_d_0 = pipe_b_311_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_d_1 = pipe_b_311_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_control_0_dataflow = mesh_7_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_control_0_propagate = mesh_7_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_control_0_shift = mesh_7_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_control_1_dataflow = mesh_7_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_control_1_propagate = mesh_7_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_control_1_shift = mesh_7_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_3_io_in_id_0 = r_567_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_3_io_in_id_1 = r_567_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_3_io_in_last_0 = r_823_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_3_io_in_last_1 = r_823_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_3_io_in_valid_0 = r_311_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_3_io_in_valid_1 = r_311_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_4_clock = clock;
  assign mesh_7_4_io_in_a_0 = r_116_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_4_io_in_a_1 = r_116_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_4_io_in_b_0 = pipe_b_71_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_b_1 = pipe_b_71_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_d_0 = pipe_b_327_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_d_1 = pipe_b_327_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_control_0_dataflow = mesh_7_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_control_0_propagate = mesh_7_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_control_0_shift = mesh_7_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_control_1_dataflow = mesh_7_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_control_1_propagate = mesh_7_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_control_1_shift = mesh_7_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_4_io_in_id_0 = r_583_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_4_io_in_id_1 = r_583_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_4_io_in_last_0 = r_839_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_4_io_in_last_1 = r_839_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_4_io_in_valid_0 = r_327_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_4_io_in_valid_1 = r_327_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_5_clock = clock;
  assign mesh_7_5_io_in_a_0 = r_117_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_5_io_in_a_1 = r_117_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_5_io_in_b_0 = pipe_b_87_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_b_1 = pipe_b_87_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_d_0 = pipe_b_343_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_d_1 = pipe_b_343_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_control_0_dataflow = mesh_7_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_control_0_propagate = mesh_7_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_control_0_shift = mesh_7_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_control_1_dataflow = mesh_7_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_control_1_propagate = mesh_7_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_control_1_shift = mesh_7_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_5_io_in_id_0 = r_599_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_5_io_in_id_1 = r_599_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_5_io_in_last_0 = r_855_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_5_io_in_last_1 = r_855_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_5_io_in_valid_0 = r_343_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_5_io_in_valid_1 = r_343_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_6_clock = clock;
  assign mesh_7_6_io_in_a_0 = r_118_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_6_io_in_a_1 = r_118_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_6_io_in_b_0 = pipe_b_103_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_b_1 = pipe_b_103_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_d_0 = pipe_b_359_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_d_1 = pipe_b_359_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_control_0_dataflow = mesh_7_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_control_0_propagate = mesh_7_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_control_0_shift = mesh_7_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_control_1_dataflow = mesh_7_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_control_1_propagate = mesh_7_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_control_1_shift = mesh_7_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_6_io_in_id_0 = r_615_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_6_io_in_id_1 = r_615_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_6_io_in_last_0 = r_871_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_6_io_in_last_1 = r_871_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_6_io_in_valid_0 = r_359_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_6_io_in_valid_1 = r_359_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_7_clock = clock;
  assign mesh_7_7_io_in_a_0 = r_119_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_7_io_in_a_1 = r_119_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_7_io_in_b_0 = pipe_b_119_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_b_1 = pipe_b_119_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_d_0 = pipe_b_375_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_d_1 = pipe_b_375_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_control_0_dataflow = mesh_7_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_control_0_propagate = mesh_7_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_control_0_shift = mesh_7_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_control_1_dataflow = mesh_7_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_control_1_propagate = mesh_7_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_control_1_shift = mesh_7_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_7_io_in_id_0 = r_631_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_7_io_in_id_1 = r_631_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_7_io_in_last_0 = r_887_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_7_io_in_last_1 = r_887_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_7_io_in_valid_0 = r_375_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_7_io_in_valid_1 = r_375_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_8_clock = clock;
  assign mesh_7_8_io_in_a_0 = r_120_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_8_io_in_a_1 = r_120_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_8_io_in_b_0 = pipe_b_135_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_b_1 = pipe_b_135_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_d_0 = pipe_b_391_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_d_1 = pipe_b_391_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_control_0_dataflow = mesh_7_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_control_0_propagate = mesh_7_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_control_0_shift = mesh_7_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_control_1_dataflow = mesh_7_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_control_1_propagate = mesh_7_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_control_1_shift = mesh_7_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_8_io_in_id_0 = r_647_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_8_io_in_id_1 = r_647_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_8_io_in_last_0 = r_903_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_8_io_in_last_1 = r_903_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_8_io_in_valid_0 = r_391_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_8_io_in_valid_1 = r_391_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_9_clock = clock;
  assign mesh_7_9_io_in_a_0 = r_121_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_9_io_in_a_1 = r_121_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_9_io_in_b_0 = pipe_b_151_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_b_1 = pipe_b_151_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_d_0 = pipe_b_407_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_d_1 = pipe_b_407_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_control_0_dataflow = mesh_7_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_control_0_propagate = mesh_7_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_control_0_shift = mesh_7_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_control_1_dataflow = mesh_7_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_control_1_propagate = mesh_7_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_control_1_shift = mesh_7_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_9_io_in_id_0 = r_663_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_9_io_in_id_1 = r_663_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_9_io_in_last_0 = r_919_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_9_io_in_last_1 = r_919_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_9_io_in_valid_0 = r_407_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_9_io_in_valid_1 = r_407_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_10_clock = clock;
  assign mesh_7_10_io_in_a_0 = r_122_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_10_io_in_a_1 = r_122_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_10_io_in_b_0 = pipe_b_167_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_b_1 = pipe_b_167_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_d_0 = pipe_b_423_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_d_1 = pipe_b_423_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_control_0_dataflow = mesh_7_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_control_0_propagate = mesh_7_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_control_0_shift = mesh_7_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_control_1_dataflow = mesh_7_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_control_1_propagate = mesh_7_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_control_1_shift = mesh_7_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_10_io_in_id_0 = r_679_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_10_io_in_id_1 = r_679_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_10_io_in_last_0 = r_935_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_10_io_in_last_1 = r_935_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_10_io_in_valid_0 = r_423_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_10_io_in_valid_1 = r_423_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_11_clock = clock;
  assign mesh_7_11_io_in_a_0 = r_123_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_11_io_in_a_1 = r_123_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_11_io_in_b_0 = pipe_b_183_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_b_1 = pipe_b_183_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_d_0 = pipe_b_439_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_d_1 = pipe_b_439_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_control_0_dataflow = mesh_7_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_control_0_propagate = mesh_7_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_control_0_shift = mesh_7_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_control_1_dataflow = mesh_7_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_control_1_propagate = mesh_7_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_control_1_shift = mesh_7_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_11_io_in_id_0 = r_695_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_11_io_in_id_1 = r_695_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_11_io_in_last_0 = r_951_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_11_io_in_last_1 = r_951_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_11_io_in_valid_0 = r_439_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_11_io_in_valid_1 = r_439_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_12_clock = clock;
  assign mesh_7_12_io_in_a_0 = r_124_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_12_io_in_a_1 = r_124_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_12_io_in_b_0 = pipe_b_199_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_b_1 = pipe_b_199_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_d_0 = pipe_b_455_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_d_1 = pipe_b_455_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_control_0_dataflow = mesh_7_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_control_0_propagate = mesh_7_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_control_0_shift = mesh_7_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_control_1_dataflow = mesh_7_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_control_1_propagate = mesh_7_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_control_1_shift = mesh_7_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_12_io_in_id_0 = r_711_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_12_io_in_id_1 = r_711_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_12_io_in_last_0 = r_967_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_12_io_in_last_1 = r_967_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_12_io_in_valid_0 = r_455_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_12_io_in_valid_1 = r_455_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_13_clock = clock;
  assign mesh_7_13_io_in_a_0 = r_125_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_13_io_in_a_1 = r_125_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_13_io_in_b_0 = pipe_b_215_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_b_1 = pipe_b_215_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_d_0 = pipe_b_471_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_d_1 = pipe_b_471_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_control_0_dataflow = mesh_7_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_control_0_propagate = mesh_7_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_control_0_shift = mesh_7_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_control_1_dataflow = mesh_7_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_control_1_propagate = mesh_7_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_control_1_shift = mesh_7_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_13_io_in_id_0 = r_727_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_13_io_in_id_1 = r_727_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_13_io_in_last_0 = r_983_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_13_io_in_last_1 = r_983_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_13_io_in_valid_0 = r_471_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_13_io_in_valid_1 = r_471_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_14_clock = clock;
  assign mesh_7_14_io_in_a_0 = r_126_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_14_io_in_a_1 = r_126_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_14_io_in_b_0 = pipe_b_231_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_b_1 = pipe_b_231_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_d_0 = pipe_b_487_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_d_1 = pipe_b_487_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_control_0_dataflow = mesh_7_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_control_0_propagate = mesh_7_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_control_0_shift = mesh_7_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_control_1_dataflow = mesh_7_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_control_1_propagate = mesh_7_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_control_1_shift = mesh_7_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_14_io_in_id_0 = r_743_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_14_io_in_id_1 = r_743_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_14_io_in_last_0 = r_999_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_14_io_in_last_1 = r_999_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_14_io_in_valid_0 = r_487_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_14_io_in_valid_1 = r_487_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_15_clock = clock;
  assign mesh_7_15_io_in_a_0 = r_127_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_15_io_in_a_1 = r_127_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_7_15_io_in_b_0 = pipe_b_247_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_b_1 = pipe_b_247_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_d_0 = pipe_b_503_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_d_1 = pipe_b_503_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_control_0_dataflow = mesh_7_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_control_0_propagate = mesh_7_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_control_0_shift = mesh_7_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_control_1_dataflow = mesh_7_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_control_1_propagate = mesh_7_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_control_1_shift = mesh_7_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_7_15_io_in_id_0 = r_759_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_15_io_in_id_1 = r_759_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_7_15_io_in_last_0 = r_1015_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_15_io_in_last_1 = r_1015_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_7_15_io_in_valid_0 = r_503_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_7_15_io_in_valid_1 = r_503_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_0_clock = clock;
  assign mesh_8_0_io_in_a_0 = r_128_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_0_io_in_a_1 = r_128_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_0_io_in_b_0 = pipe_b_8_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_b_1 = pipe_b_8_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_d_0 = pipe_b_264_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_d_1 = pipe_b_264_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_control_0_dataflow = mesh_8_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_control_0_propagate = mesh_8_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_control_0_shift = mesh_8_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_control_1_dataflow = mesh_8_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_control_1_propagate = mesh_8_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_control_1_shift = mesh_8_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_0_io_in_id_0 = r_520_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_0_io_in_id_1 = r_520_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_0_io_in_last_0 = r_776_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_0_io_in_last_1 = r_776_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_0_io_in_valid_0 = r_264_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_0_io_in_valid_1 = r_264_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_1_clock = clock;
  assign mesh_8_1_io_in_a_0 = r_129_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_1_io_in_a_1 = r_129_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_1_io_in_b_0 = pipe_b_24_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_b_1 = pipe_b_24_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_d_0 = pipe_b_280_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_d_1 = pipe_b_280_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_control_0_dataflow = mesh_8_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_control_0_propagate = mesh_8_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_control_0_shift = mesh_8_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_control_1_dataflow = mesh_8_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_control_1_propagate = mesh_8_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_control_1_shift = mesh_8_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_1_io_in_id_0 = r_536_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_1_io_in_id_1 = r_536_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_1_io_in_last_0 = r_792_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_1_io_in_last_1 = r_792_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_1_io_in_valid_0 = r_280_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_1_io_in_valid_1 = r_280_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_2_clock = clock;
  assign mesh_8_2_io_in_a_0 = r_130_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_2_io_in_a_1 = r_130_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_2_io_in_b_0 = pipe_b_40_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_b_1 = pipe_b_40_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_d_0 = pipe_b_296_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_d_1 = pipe_b_296_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_control_0_dataflow = mesh_8_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_control_0_propagate = mesh_8_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_control_0_shift = mesh_8_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_control_1_dataflow = mesh_8_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_control_1_propagate = mesh_8_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_control_1_shift = mesh_8_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_2_io_in_id_0 = r_552_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_2_io_in_id_1 = r_552_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_2_io_in_last_0 = r_808_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_2_io_in_last_1 = r_808_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_2_io_in_valid_0 = r_296_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_2_io_in_valid_1 = r_296_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_3_clock = clock;
  assign mesh_8_3_io_in_a_0 = r_131_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_3_io_in_a_1 = r_131_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_3_io_in_b_0 = pipe_b_56_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_b_1 = pipe_b_56_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_d_0 = pipe_b_312_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_d_1 = pipe_b_312_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_control_0_dataflow = mesh_8_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_control_0_propagate = mesh_8_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_control_0_shift = mesh_8_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_control_1_dataflow = mesh_8_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_control_1_propagate = mesh_8_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_control_1_shift = mesh_8_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_3_io_in_id_0 = r_568_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_3_io_in_id_1 = r_568_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_3_io_in_last_0 = r_824_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_3_io_in_last_1 = r_824_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_3_io_in_valid_0 = r_312_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_3_io_in_valid_1 = r_312_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_4_clock = clock;
  assign mesh_8_4_io_in_a_0 = r_132_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_4_io_in_a_1 = r_132_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_4_io_in_b_0 = pipe_b_72_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_b_1 = pipe_b_72_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_d_0 = pipe_b_328_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_d_1 = pipe_b_328_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_control_0_dataflow = mesh_8_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_control_0_propagate = mesh_8_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_control_0_shift = mesh_8_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_control_1_dataflow = mesh_8_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_control_1_propagate = mesh_8_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_control_1_shift = mesh_8_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_4_io_in_id_0 = r_584_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_4_io_in_id_1 = r_584_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_4_io_in_last_0 = r_840_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_4_io_in_last_1 = r_840_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_4_io_in_valid_0 = r_328_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_4_io_in_valid_1 = r_328_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_5_clock = clock;
  assign mesh_8_5_io_in_a_0 = r_133_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_5_io_in_a_1 = r_133_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_5_io_in_b_0 = pipe_b_88_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_b_1 = pipe_b_88_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_d_0 = pipe_b_344_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_d_1 = pipe_b_344_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_control_0_dataflow = mesh_8_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_control_0_propagate = mesh_8_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_control_0_shift = mesh_8_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_control_1_dataflow = mesh_8_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_control_1_propagate = mesh_8_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_control_1_shift = mesh_8_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_5_io_in_id_0 = r_600_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_5_io_in_id_1 = r_600_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_5_io_in_last_0 = r_856_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_5_io_in_last_1 = r_856_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_5_io_in_valid_0 = r_344_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_5_io_in_valid_1 = r_344_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_6_clock = clock;
  assign mesh_8_6_io_in_a_0 = r_134_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_6_io_in_a_1 = r_134_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_6_io_in_b_0 = pipe_b_104_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_b_1 = pipe_b_104_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_d_0 = pipe_b_360_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_d_1 = pipe_b_360_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_control_0_dataflow = mesh_8_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_control_0_propagate = mesh_8_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_control_0_shift = mesh_8_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_control_1_dataflow = mesh_8_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_control_1_propagate = mesh_8_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_control_1_shift = mesh_8_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_6_io_in_id_0 = r_616_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_6_io_in_id_1 = r_616_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_6_io_in_last_0 = r_872_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_6_io_in_last_1 = r_872_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_6_io_in_valid_0 = r_360_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_6_io_in_valid_1 = r_360_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_7_clock = clock;
  assign mesh_8_7_io_in_a_0 = r_135_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_7_io_in_a_1 = r_135_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_7_io_in_b_0 = pipe_b_120_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_b_1 = pipe_b_120_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_d_0 = pipe_b_376_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_d_1 = pipe_b_376_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_control_0_dataflow = mesh_8_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_control_0_propagate = mesh_8_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_control_0_shift = mesh_8_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_control_1_dataflow = mesh_8_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_control_1_propagate = mesh_8_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_control_1_shift = mesh_8_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_7_io_in_id_0 = r_632_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_7_io_in_id_1 = r_632_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_7_io_in_last_0 = r_888_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_7_io_in_last_1 = r_888_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_7_io_in_valid_0 = r_376_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_7_io_in_valid_1 = r_376_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_8_clock = clock;
  assign mesh_8_8_io_in_a_0 = r_136_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_8_io_in_a_1 = r_136_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_8_io_in_b_0 = pipe_b_136_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_b_1 = pipe_b_136_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_d_0 = pipe_b_392_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_d_1 = pipe_b_392_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_control_0_dataflow = mesh_8_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_control_0_propagate = mesh_8_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_control_0_shift = mesh_8_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_control_1_dataflow = mesh_8_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_control_1_propagate = mesh_8_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_control_1_shift = mesh_8_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_8_io_in_id_0 = r_648_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_8_io_in_id_1 = r_648_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_8_io_in_last_0 = r_904_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_8_io_in_last_1 = r_904_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_8_io_in_valid_0 = r_392_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_8_io_in_valid_1 = r_392_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_9_clock = clock;
  assign mesh_8_9_io_in_a_0 = r_137_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_9_io_in_a_1 = r_137_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_9_io_in_b_0 = pipe_b_152_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_b_1 = pipe_b_152_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_d_0 = pipe_b_408_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_d_1 = pipe_b_408_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_control_0_dataflow = mesh_8_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_control_0_propagate = mesh_8_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_control_0_shift = mesh_8_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_control_1_dataflow = mesh_8_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_control_1_propagate = mesh_8_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_control_1_shift = mesh_8_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_9_io_in_id_0 = r_664_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_9_io_in_id_1 = r_664_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_9_io_in_last_0 = r_920_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_9_io_in_last_1 = r_920_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_9_io_in_valid_0 = r_408_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_9_io_in_valid_1 = r_408_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_10_clock = clock;
  assign mesh_8_10_io_in_a_0 = r_138_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_10_io_in_a_1 = r_138_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_10_io_in_b_0 = pipe_b_168_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_b_1 = pipe_b_168_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_d_0 = pipe_b_424_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_d_1 = pipe_b_424_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_control_0_dataflow = mesh_8_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_control_0_propagate = mesh_8_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_control_0_shift = mesh_8_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_control_1_dataflow = mesh_8_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_control_1_propagate = mesh_8_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_control_1_shift = mesh_8_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_10_io_in_id_0 = r_680_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_10_io_in_id_1 = r_680_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_10_io_in_last_0 = r_936_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_10_io_in_last_1 = r_936_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_10_io_in_valid_0 = r_424_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_10_io_in_valid_1 = r_424_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_11_clock = clock;
  assign mesh_8_11_io_in_a_0 = r_139_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_11_io_in_a_1 = r_139_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_11_io_in_b_0 = pipe_b_184_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_b_1 = pipe_b_184_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_d_0 = pipe_b_440_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_d_1 = pipe_b_440_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_control_0_dataflow = mesh_8_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_control_0_propagate = mesh_8_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_control_0_shift = mesh_8_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_control_1_dataflow = mesh_8_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_control_1_propagate = mesh_8_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_control_1_shift = mesh_8_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_11_io_in_id_0 = r_696_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_11_io_in_id_1 = r_696_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_11_io_in_last_0 = r_952_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_11_io_in_last_1 = r_952_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_11_io_in_valid_0 = r_440_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_11_io_in_valid_1 = r_440_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_12_clock = clock;
  assign mesh_8_12_io_in_a_0 = r_140_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_12_io_in_a_1 = r_140_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_12_io_in_b_0 = pipe_b_200_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_b_1 = pipe_b_200_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_d_0 = pipe_b_456_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_d_1 = pipe_b_456_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_control_0_dataflow = mesh_8_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_control_0_propagate = mesh_8_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_control_0_shift = mesh_8_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_control_1_dataflow = mesh_8_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_control_1_propagate = mesh_8_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_control_1_shift = mesh_8_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_12_io_in_id_0 = r_712_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_12_io_in_id_1 = r_712_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_12_io_in_last_0 = r_968_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_12_io_in_last_1 = r_968_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_12_io_in_valid_0 = r_456_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_12_io_in_valid_1 = r_456_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_13_clock = clock;
  assign mesh_8_13_io_in_a_0 = r_141_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_13_io_in_a_1 = r_141_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_13_io_in_b_0 = pipe_b_216_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_b_1 = pipe_b_216_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_d_0 = pipe_b_472_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_d_1 = pipe_b_472_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_control_0_dataflow = mesh_8_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_control_0_propagate = mesh_8_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_control_0_shift = mesh_8_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_control_1_dataflow = mesh_8_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_control_1_propagate = mesh_8_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_control_1_shift = mesh_8_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_13_io_in_id_0 = r_728_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_13_io_in_id_1 = r_728_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_13_io_in_last_0 = r_984_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_13_io_in_last_1 = r_984_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_13_io_in_valid_0 = r_472_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_13_io_in_valid_1 = r_472_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_14_clock = clock;
  assign mesh_8_14_io_in_a_0 = r_142_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_14_io_in_a_1 = r_142_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_14_io_in_b_0 = pipe_b_232_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_b_1 = pipe_b_232_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_d_0 = pipe_b_488_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_d_1 = pipe_b_488_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_control_0_dataflow = mesh_8_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_control_0_propagate = mesh_8_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_control_0_shift = mesh_8_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_control_1_dataflow = mesh_8_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_control_1_propagate = mesh_8_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_control_1_shift = mesh_8_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_14_io_in_id_0 = r_744_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_14_io_in_id_1 = r_744_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_14_io_in_last_0 = r_1000_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_14_io_in_last_1 = r_1000_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_14_io_in_valid_0 = r_488_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_14_io_in_valid_1 = r_488_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_15_clock = clock;
  assign mesh_8_15_io_in_a_0 = r_143_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_15_io_in_a_1 = r_143_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_8_15_io_in_b_0 = pipe_b_248_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_b_1 = pipe_b_248_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_d_0 = pipe_b_504_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_d_1 = pipe_b_504_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_control_0_dataflow = mesh_8_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_control_0_propagate = mesh_8_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_control_0_shift = mesh_8_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_control_1_dataflow = mesh_8_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_control_1_propagate = mesh_8_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_control_1_shift = mesh_8_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_8_15_io_in_id_0 = r_760_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_15_io_in_id_1 = r_760_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_8_15_io_in_last_0 = r_1016_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_15_io_in_last_1 = r_1016_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_8_15_io_in_valid_0 = r_504_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_8_15_io_in_valid_1 = r_504_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_0_clock = clock;
  assign mesh_9_0_io_in_a_0 = r_144_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_0_io_in_a_1 = r_144_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_0_io_in_b_0 = pipe_b_9_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_b_1 = pipe_b_9_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_d_0 = pipe_b_265_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_d_1 = pipe_b_265_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_control_0_dataflow = mesh_9_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_control_0_propagate = mesh_9_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_control_0_shift = mesh_9_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_control_1_dataflow = mesh_9_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_control_1_propagate = mesh_9_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_control_1_shift = mesh_9_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_0_io_in_id_0 = r_521_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_0_io_in_id_1 = r_521_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_0_io_in_last_0 = r_777_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_0_io_in_last_1 = r_777_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_0_io_in_valid_0 = r_265_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_0_io_in_valid_1 = r_265_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_1_clock = clock;
  assign mesh_9_1_io_in_a_0 = r_145_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_1_io_in_a_1 = r_145_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_1_io_in_b_0 = pipe_b_25_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_b_1 = pipe_b_25_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_d_0 = pipe_b_281_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_d_1 = pipe_b_281_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_control_0_dataflow = mesh_9_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_control_0_propagate = mesh_9_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_control_0_shift = mesh_9_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_control_1_dataflow = mesh_9_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_control_1_propagate = mesh_9_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_control_1_shift = mesh_9_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_1_io_in_id_0 = r_537_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_1_io_in_id_1 = r_537_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_1_io_in_last_0 = r_793_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_1_io_in_last_1 = r_793_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_1_io_in_valid_0 = r_281_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_1_io_in_valid_1 = r_281_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_2_clock = clock;
  assign mesh_9_2_io_in_a_0 = r_146_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_2_io_in_a_1 = r_146_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_2_io_in_b_0 = pipe_b_41_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_b_1 = pipe_b_41_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_d_0 = pipe_b_297_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_d_1 = pipe_b_297_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_control_0_dataflow = mesh_9_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_control_0_propagate = mesh_9_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_control_0_shift = mesh_9_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_control_1_dataflow = mesh_9_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_control_1_propagate = mesh_9_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_control_1_shift = mesh_9_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_2_io_in_id_0 = r_553_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_2_io_in_id_1 = r_553_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_2_io_in_last_0 = r_809_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_2_io_in_last_1 = r_809_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_2_io_in_valid_0 = r_297_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_2_io_in_valid_1 = r_297_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_3_clock = clock;
  assign mesh_9_3_io_in_a_0 = r_147_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_3_io_in_a_1 = r_147_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_3_io_in_b_0 = pipe_b_57_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_b_1 = pipe_b_57_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_d_0 = pipe_b_313_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_d_1 = pipe_b_313_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_control_0_dataflow = mesh_9_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_control_0_propagate = mesh_9_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_control_0_shift = mesh_9_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_control_1_dataflow = mesh_9_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_control_1_propagate = mesh_9_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_control_1_shift = mesh_9_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_3_io_in_id_0 = r_569_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_3_io_in_id_1 = r_569_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_3_io_in_last_0 = r_825_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_3_io_in_last_1 = r_825_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_3_io_in_valid_0 = r_313_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_3_io_in_valid_1 = r_313_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_4_clock = clock;
  assign mesh_9_4_io_in_a_0 = r_148_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_4_io_in_a_1 = r_148_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_4_io_in_b_0 = pipe_b_73_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_b_1 = pipe_b_73_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_d_0 = pipe_b_329_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_d_1 = pipe_b_329_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_control_0_dataflow = mesh_9_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_control_0_propagate = mesh_9_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_control_0_shift = mesh_9_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_control_1_dataflow = mesh_9_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_control_1_propagate = mesh_9_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_control_1_shift = mesh_9_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_4_io_in_id_0 = r_585_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_4_io_in_id_1 = r_585_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_4_io_in_last_0 = r_841_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_4_io_in_last_1 = r_841_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_4_io_in_valid_0 = r_329_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_4_io_in_valid_1 = r_329_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_5_clock = clock;
  assign mesh_9_5_io_in_a_0 = r_149_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_5_io_in_a_1 = r_149_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_5_io_in_b_0 = pipe_b_89_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_b_1 = pipe_b_89_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_d_0 = pipe_b_345_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_d_1 = pipe_b_345_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_control_0_dataflow = mesh_9_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_control_0_propagate = mesh_9_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_control_0_shift = mesh_9_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_control_1_dataflow = mesh_9_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_control_1_propagate = mesh_9_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_control_1_shift = mesh_9_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_5_io_in_id_0 = r_601_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_5_io_in_id_1 = r_601_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_5_io_in_last_0 = r_857_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_5_io_in_last_1 = r_857_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_5_io_in_valid_0 = r_345_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_5_io_in_valid_1 = r_345_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_6_clock = clock;
  assign mesh_9_6_io_in_a_0 = r_150_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_6_io_in_a_1 = r_150_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_6_io_in_b_0 = pipe_b_105_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_b_1 = pipe_b_105_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_d_0 = pipe_b_361_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_d_1 = pipe_b_361_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_control_0_dataflow = mesh_9_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_control_0_propagate = mesh_9_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_control_0_shift = mesh_9_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_control_1_dataflow = mesh_9_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_control_1_propagate = mesh_9_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_control_1_shift = mesh_9_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_6_io_in_id_0 = r_617_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_6_io_in_id_1 = r_617_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_6_io_in_last_0 = r_873_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_6_io_in_last_1 = r_873_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_6_io_in_valid_0 = r_361_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_6_io_in_valid_1 = r_361_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_7_clock = clock;
  assign mesh_9_7_io_in_a_0 = r_151_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_7_io_in_a_1 = r_151_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_7_io_in_b_0 = pipe_b_121_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_b_1 = pipe_b_121_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_d_0 = pipe_b_377_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_d_1 = pipe_b_377_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_control_0_dataflow = mesh_9_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_control_0_propagate = mesh_9_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_control_0_shift = mesh_9_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_control_1_dataflow = mesh_9_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_control_1_propagate = mesh_9_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_control_1_shift = mesh_9_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_7_io_in_id_0 = r_633_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_7_io_in_id_1 = r_633_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_7_io_in_last_0 = r_889_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_7_io_in_last_1 = r_889_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_7_io_in_valid_0 = r_377_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_7_io_in_valid_1 = r_377_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_8_clock = clock;
  assign mesh_9_8_io_in_a_0 = r_152_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_8_io_in_a_1 = r_152_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_8_io_in_b_0 = pipe_b_137_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_b_1 = pipe_b_137_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_d_0 = pipe_b_393_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_d_1 = pipe_b_393_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_control_0_dataflow = mesh_9_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_control_0_propagate = mesh_9_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_control_0_shift = mesh_9_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_control_1_dataflow = mesh_9_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_control_1_propagate = mesh_9_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_control_1_shift = mesh_9_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_8_io_in_id_0 = r_649_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_8_io_in_id_1 = r_649_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_8_io_in_last_0 = r_905_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_8_io_in_last_1 = r_905_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_8_io_in_valid_0 = r_393_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_8_io_in_valid_1 = r_393_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_9_clock = clock;
  assign mesh_9_9_io_in_a_0 = r_153_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_9_io_in_a_1 = r_153_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_9_io_in_b_0 = pipe_b_153_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_b_1 = pipe_b_153_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_d_0 = pipe_b_409_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_d_1 = pipe_b_409_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_control_0_dataflow = mesh_9_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_control_0_propagate = mesh_9_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_control_0_shift = mesh_9_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_control_1_dataflow = mesh_9_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_control_1_propagate = mesh_9_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_control_1_shift = mesh_9_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_9_io_in_id_0 = r_665_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_9_io_in_id_1 = r_665_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_9_io_in_last_0 = r_921_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_9_io_in_last_1 = r_921_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_9_io_in_valid_0 = r_409_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_9_io_in_valid_1 = r_409_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_10_clock = clock;
  assign mesh_9_10_io_in_a_0 = r_154_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_10_io_in_a_1 = r_154_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_10_io_in_b_0 = pipe_b_169_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_b_1 = pipe_b_169_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_d_0 = pipe_b_425_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_d_1 = pipe_b_425_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_control_0_dataflow = mesh_9_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_control_0_propagate = mesh_9_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_control_0_shift = mesh_9_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_control_1_dataflow = mesh_9_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_control_1_propagate = mesh_9_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_control_1_shift = mesh_9_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_10_io_in_id_0 = r_681_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_10_io_in_id_1 = r_681_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_10_io_in_last_0 = r_937_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_10_io_in_last_1 = r_937_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_10_io_in_valid_0 = r_425_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_10_io_in_valid_1 = r_425_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_11_clock = clock;
  assign mesh_9_11_io_in_a_0 = r_155_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_11_io_in_a_1 = r_155_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_11_io_in_b_0 = pipe_b_185_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_b_1 = pipe_b_185_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_d_0 = pipe_b_441_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_d_1 = pipe_b_441_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_control_0_dataflow = mesh_9_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_control_0_propagate = mesh_9_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_control_0_shift = mesh_9_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_control_1_dataflow = mesh_9_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_control_1_propagate = mesh_9_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_control_1_shift = mesh_9_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_11_io_in_id_0 = r_697_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_11_io_in_id_1 = r_697_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_11_io_in_last_0 = r_953_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_11_io_in_last_1 = r_953_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_11_io_in_valid_0 = r_441_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_11_io_in_valid_1 = r_441_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_12_clock = clock;
  assign mesh_9_12_io_in_a_0 = r_156_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_12_io_in_a_1 = r_156_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_12_io_in_b_0 = pipe_b_201_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_b_1 = pipe_b_201_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_d_0 = pipe_b_457_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_d_1 = pipe_b_457_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_control_0_dataflow = mesh_9_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_control_0_propagate = mesh_9_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_control_0_shift = mesh_9_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_control_1_dataflow = mesh_9_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_control_1_propagate = mesh_9_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_control_1_shift = mesh_9_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_12_io_in_id_0 = r_713_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_12_io_in_id_1 = r_713_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_12_io_in_last_0 = r_969_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_12_io_in_last_1 = r_969_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_12_io_in_valid_0 = r_457_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_12_io_in_valid_1 = r_457_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_13_clock = clock;
  assign mesh_9_13_io_in_a_0 = r_157_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_13_io_in_a_1 = r_157_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_13_io_in_b_0 = pipe_b_217_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_b_1 = pipe_b_217_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_d_0 = pipe_b_473_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_d_1 = pipe_b_473_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_control_0_dataflow = mesh_9_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_control_0_propagate = mesh_9_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_control_0_shift = mesh_9_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_control_1_dataflow = mesh_9_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_control_1_propagate = mesh_9_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_control_1_shift = mesh_9_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_13_io_in_id_0 = r_729_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_13_io_in_id_1 = r_729_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_13_io_in_last_0 = r_985_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_13_io_in_last_1 = r_985_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_13_io_in_valid_0 = r_473_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_13_io_in_valid_1 = r_473_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_14_clock = clock;
  assign mesh_9_14_io_in_a_0 = r_158_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_14_io_in_a_1 = r_158_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_14_io_in_b_0 = pipe_b_233_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_b_1 = pipe_b_233_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_d_0 = pipe_b_489_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_d_1 = pipe_b_489_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_control_0_dataflow = mesh_9_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_control_0_propagate = mesh_9_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_control_0_shift = mesh_9_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_control_1_dataflow = mesh_9_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_control_1_propagate = mesh_9_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_control_1_shift = mesh_9_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_14_io_in_id_0 = r_745_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_14_io_in_id_1 = r_745_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_14_io_in_last_0 = r_1001_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_14_io_in_last_1 = r_1001_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_14_io_in_valid_0 = r_489_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_14_io_in_valid_1 = r_489_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_15_clock = clock;
  assign mesh_9_15_io_in_a_0 = r_159_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_15_io_in_a_1 = r_159_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_9_15_io_in_b_0 = pipe_b_249_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_b_1 = pipe_b_249_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_d_0 = pipe_b_505_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_d_1 = pipe_b_505_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_control_0_dataflow = mesh_9_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_control_0_propagate = mesh_9_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_control_0_shift = mesh_9_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_control_1_dataflow = mesh_9_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_control_1_propagate = mesh_9_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_control_1_shift = mesh_9_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_9_15_io_in_id_0 = r_761_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_15_io_in_id_1 = r_761_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_9_15_io_in_last_0 = r_1017_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_15_io_in_last_1 = r_1017_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_9_15_io_in_valid_0 = r_505_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_9_15_io_in_valid_1 = r_505_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_0_clock = clock;
  assign mesh_10_0_io_in_a_0 = r_160_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_0_io_in_a_1 = r_160_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_0_io_in_b_0 = pipe_b_10_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_b_1 = pipe_b_10_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_d_0 = pipe_b_266_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_d_1 = pipe_b_266_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_control_0_dataflow = mesh_10_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_control_0_propagate = mesh_10_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_control_0_shift = mesh_10_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_control_1_dataflow = mesh_10_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_control_1_propagate = mesh_10_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_control_1_shift = mesh_10_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_0_io_in_id_0 = r_522_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_0_io_in_id_1 = r_522_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_0_io_in_last_0 = r_778_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_0_io_in_last_1 = r_778_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_0_io_in_valid_0 = r_266_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_0_io_in_valid_1 = r_266_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_1_clock = clock;
  assign mesh_10_1_io_in_a_0 = r_161_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_1_io_in_a_1 = r_161_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_1_io_in_b_0 = pipe_b_26_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_b_1 = pipe_b_26_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_d_0 = pipe_b_282_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_d_1 = pipe_b_282_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_control_0_dataflow = mesh_10_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_control_0_propagate = mesh_10_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_control_0_shift = mesh_10_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_control_1_dataflow = mesh_10_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_control_1_propagate = mesh_10_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_control_1_shift = mesh_10_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_1_io_in_id_0 = r_538_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_1_io_in_id_1 = r_538_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_1_io_in_last_0 = r_794_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_1_io_in_last_1 = r_794_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_1_io_in_valid_0 = r_282_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_1_io_in_valid_1 = r_282_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_2_clock = clock;
  assign mesh_10_2_io_in_a_0 = r_162_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_2_io_in_a_1 = r_162_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_2_io_in_b_0 = pipe_b_42_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_b_1 = pipe_b_42_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_d_0 = pipe_b_298_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_d_1 = pipe_b_298_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_control_0_dataflow = mesh_10_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_control_0_propagate = mesh_10_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_control_0_shift = mesh_10_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_control_1_dataflow = mesh_10_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_control_1_propagate = mesh_10_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_control_1_shift = mesh_10_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_2_io_in_id_0 = r_554_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_2_io_in_id_1 = r_554_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_2_io_in_last_0 = r_810_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_2_io_in_last_1 = r_810_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_2_io_in_valid_0 = r_298_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_2_io_in_valid_1 = r_298_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_3_clock = clock;
  assign mesh_10_3_io_in_a_0 = r_163_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_3_io_in_a_1 = r_163_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_3_io_in_b_0 = pipe_b_58_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_b_1 = pipe_b_58_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_d_0 = pipe_b_314_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_d_1 = pipe_b_314_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_control_0_dataflow = mesh_10_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_control_0_propagate = mesh_10_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_control_0_shift = mesh_10_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_control_1_dataflow = mesh_10_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_control_1_propagate = mesh_10_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_control_1_shift = mesh_10_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_3_io_in_id_0 = r_570_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_3_io_in_id_1 = r_570_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_3_io_in_last_0 = r_826_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_3_io_in_last_1 = r_826_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_3_io_in_valid_0 = r_314_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_3_io_in_valid_1 = r_314_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_4_clock = clock;
  assign mesh_10_4_io_in_a_0 = r_164_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_4_io_in_a_1 = r_164_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_4_io_in_b_0 = pipe_b_74_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_b_1 = pipe_b_74_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_d_0 = pipe_b_330_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_d_1 = pipe_b_330_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_control_0_dataflow = mesh_10_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_control_0_propagate = mesh_10_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_control_0_shift = mesh_10_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_control_1_dataflow = mesh_10_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_control_1_propagate = mesh_10_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_control_1_shift = mesh_10_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_4_io_in_id_0 = r_586_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_4_io_in_id_1 = r_586_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_4_io_in_last_0 = r_842_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_4_io_in_last_1 = r_842_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_4_io_in_valid_0 = r_330_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_4_io_in_valid_1 = r_330_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_5_clock = clock;
  assign mesh_10_5_io_in_a_0 = r_165_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_5_io_in_a_1 = r_165_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_5_io_in_b_0 = pipe_b_90_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_b_1 = pipe_b_90_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_d_0 = pipe_b_346_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_d_1 = pipe_b_346_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_control_0_dataflow = mesh_10_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_control_0_propagate = mesh_10_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_control_0_shift = mesh_10_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_control_1_dataflow = mesh_10_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_control_1_propagate = mesh_10_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_control_1_shift = mesh_10_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_5_io_in_id_0 = r_602_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_5_io_in_id_1 = r_602_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_5_io_in_last_0 = r_858_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_5_io_in_last_1 = r_858_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_5_io_in_valid_0 = r_346_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_5_io_in_valid_1 = r_346_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_6_clock = clock;
  assign mesh_10_6_io_in_a_0 = r_166_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_6_io_in_a_1 = r_166_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_6_io_in_b_0 = pipe_b_106_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_b_1 = pipe_b_106_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_d_0 = pipe_b_362_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_d_1 = pipe_b_362_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_control_0_dataflow = mesh_10_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_control_0_propagate = mesh_10_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_control_0_shift = mesh_10_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_control_1_dataflow = mesh_10_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_control_1_propagate = mesh_10_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_control_1_shift = mesh_10_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_6_io_in_id_0 = r_618_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_6_io_in_id_1 = r_618_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_6_io_in_last_0 = r_874_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_6_io_in_last_1 = r_874_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_6_io_in_valid_0 = r_362_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_6_io_in_valid_1 = r_362_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_7_clock = clock;
  assign mesh_10_7_io_in_a_0 = r_167_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_7_io_in_a_1 = r_167_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_7_io_in_b_0 = pipe_b_122_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_b_1 = pipe_b_122_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_d_0 = pipe_b_378_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_d_1 = pipe_b_378_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_control_0_dataflow = mesh_10_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_control_0_propagate = mesh_10_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_control_0_shift = mesh_10_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_control_1_dataflow = mesh_10_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_control_1_propagate = mesh_10_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_control_1_shift = mesh_10_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_7_io_in_id_0 = r_634_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_7_io_in_id_1 = r_634_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_7_io_in_last_0 = r_890_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_7_io_in_last_1 = r_890_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_7_io_in_valid_0 = r_378_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_7_io_in_valid_1 = r_378_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_8_clock = clock;
  assign mesh_10_8_io_in_a_0 = r_168_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_8_io_in_a_1 = r_168_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_8_io_in_b_0 = pipe_b_138_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_b_1 = pipe_b_138_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_d_0 = pipe_b_394_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_d_1 = pipe_b_394_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_control_0_dataflow = mesh_10_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_control_0_propagate = mesh_10_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_control_0_shift = mesh_10_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_control_1_dataflow = mesh_10_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_control_1_propagate = mesh_10_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_control_1_shift = mesh_10_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_8_io_in_id_0 = r_650_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_8_io_in_id_1 = r_650_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_8_io_in_last_0 = r_906_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_8_io_in_last_1 = r_906_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_8_io_in_valid_0 = r_394_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_8_io_in_valid_1 = r_394_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_9_clock = clock;
  assign mesh_10_9_io_in_a_0 = r_169_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_9_io_in_a_1 = r_169_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_9_io_in_b_0 = pipe_b_154_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_b_1 = pipe_b_154_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_d_0 = pipe_b_410_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_d_1 = pipe_b_410_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_control_0_dataflow = mesh_10_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_control_0_propagate = mesh_10_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_control_0_shift = mesh_10_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_control_1_dataflow = mesh_10_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_control_1_propagate = mesh_10_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_control_1_shift = mesh_10_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_9_io_in_id_0 = r_666_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_9_io_in_id_1 = r_666_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_9_io_in_last_0 = r_922_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_9_io_in_last_1 = r_922_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_9_io_in_valid_0 = r_410_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_9_io_in_valid_1 = r_410_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_10_clock = clock;
  assign mesh_10_10_io_in_a_0 = r_170_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_10_io_in_a_1 = r_170_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_10_io_in_b_0 = pipe_b_170_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_b_1 = pipe_b_170_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_d_0 = pipe_b_426_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_d_1 = pipe_b_426_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_control_0_dataflow = mesh_10_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_control_0_propagate = mesh_10_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_control_0_shift = mesh_10_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_control_1_dataflow = mesh_10_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_control_1_propagate = mesh_10_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_control_1_shift = mesh_10_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_10_io_in_id_0 = r_682_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_10_io_in_id_1 = r_682_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_10_io_in_last_0 = r_938_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_10_io_in_last_1 = r_938_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_10_io_in_valid_0 = r_426_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_10_io_in_valid_1 = r_426_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_11_clock = clock;
  assign mesh_10_11_io_in_a_0 = r_171_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_11_io_in_a_1 = r_171_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_11_io_in_b_0 = pipe_b_186_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_b_1 = pipe_b_186_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_d_0 = pipe_b_442_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_d_1 = pipe_b_442_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_control_0_dataflow = mesh_10_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_control_0_propagate = mesh_10_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_control_0_shift = mesh_10_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_control_1_dataflow = mesh_10_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_control_1_propagate = mesh_10_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_control_1_shift = mesh_10_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_11_io_in_id_0 = r_698_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_11_io_in_id_1 = r_698_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_11_io_in_last_0 = r_954_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_11_io_in_last_1 = r_954_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_11_io_in_valid_0 = r_442_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_11_io_in_valid_1 = r_442_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_12_clock = clock;
  assign mesh_10_12_io_in_a_0 = r_172_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_12_io_in_a_1 = r_172_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_12_io_in_b_0 = pipe_b_202_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_b_1 = pipe_b_202_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_d_0 = pipe_b_458_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_d_1 = pipe_b_458_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_control_0_dataflow = mesh_10_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_control_0_propagate = mesh_10_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_control_0_shift = mesh_10_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_control_1_dataflow = mesh_10_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_control_1_propagate = mesh_10_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_control_1_shift = mesh_10_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_12_io_in_id_0 = r_714_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_12_io_in_id_1 = r_714_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_12_io_in_last_0 = r_970_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_12_io_in_last_1 = r_970_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_12_io_in_valid_0 = r_458_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_12_io_in_valid_1 = r_458_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_13_clock = clock;
  assign mesh_10_13_io_in_a_0 = r_173_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_13_io_in_a_1 = r_173_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_13_io_in_b_0 = pipe_b_218_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_b_1 = pipe_b_218_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_d_0 = pipe_b_474_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_d_1 = pipe_b_474_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_control_0_dataflow = mesh_10_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_control_0_propagate = mesh_10_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_control_0_shift = mesh_10_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_control_1_dataflow = mesh_10_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_control_1_propagate = mesh_10_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_control_1_shift = mesh_10_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_13_io_in_id_0 = r_730_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_13_io_in_id_1 = r_730_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_13_io_in_last_0 = r_986_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_13_io_in_last_1 = r_986_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_13_io_in_valid_0 = r_474_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_13_io_in_valid_1 = r_474_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_14_clock = clock;
  assign mesh_10_14_io_in_a_0 = r_174_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_14_io_in_a_1 = r_174_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_14_io_in_b_0 = pipe_b_234_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_b_1 = pipe_b_234_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_d_0 = pipe_b_490_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_d_1 = pipe_b_490_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_control_0_dataflow = mesh_10_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_control_0_propagate = mesh_10_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_control_0_shift = mesh_10_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_control_1_dataflow = mesh_10_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_control_1_propagate = mesh_10_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_control_1_shift = mesh_10_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_14_io_in_id_0 = r_746_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_14_io_in_id_1 = r_746_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_14_io_in_last_0 = r_1002_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_14_io_in_last_1 = r_1002_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_14_io_in_valid_0 = r_490_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_14_io_in_valid_1 = r_490_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_15_clock = clock;
  assign mesh_10_15_io_in_a_0 = r_175_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_15_io_in_a_1 = r_175_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_10_15_io_in_b_0 = pipe_b_250_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_b_1 = pipe_b_250_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_d_0 = pipe_b_506_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_d_1 = pipe_b_506_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_control_0_dataflow = mesh_10_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_control_0_propagate = mesh_10_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_control_0_shift = mesh_10_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_control_1_dataflow = mesh_10_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_control_1_propagate = mesh_10_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_control_1_shift = mesh_10_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_10_15_io_in_id_0 = r_762_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_15_io_in_id_1 = r_762_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_10_15_io_in_last_0 = r_1018_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_15_io_in_last_1 = r_1018_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_10_15_io_in_valid_0 = r_506_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_10_15_io_in_valid_1 = r_506_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_0_clock = clock;
  assign mesh_11_0_io_in_a_0 = r_176_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_0_io_in_a_1 = r_176_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_0_io_in_b_0 = pipe_b_11_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_b_1 = pipe_b_11_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_d_0 = pipe_b_267_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_d_1 = pipe_b_267_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_control_0_dataflow = mesh_11_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_control_0_propagate = mesh_11_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_control_0_shift = mesh_11_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_control_1_dataflow = mesh_11_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_control_1_propagate = mesh_11_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_control_1_shift = mesh_11_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_0_io_in_id_0 = r_523_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_0_io_in_id_1 = r_523_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_0_io_in_last_0 = r_779_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_0_io_in_last_1 = r_779_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_0_io_in_valid_0 = r_267_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_0_io_in_valid_1 = r_267_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_1_clock = clock;
  assign mesh_11_1_io_in_a_0 = r_177_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_1_io_in_a_1 = r_177_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_1_io_in_b_0 = pipe_b_27_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_b_1 = pipe_b_27_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_d_0 = pipe_b_283_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_d_1 = pipe_b_283_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_control_0_dataflow = mesh_11_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_control_0_propagate = mesh_11_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_control_0_shift = mesh_11_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_control_1_dataflow = mesh_11_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_control_1_propagate = mesh_11_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_control_1_shift = mesh_11_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_1_io_in_id_0 = r_539_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_1_io_in_id_1 = r_539_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_1_io_in_last_0 = r_795_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_1_io_in_last_1 = r_795_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_1_io_in_valid_0 = r_283_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_1_io_in_valid_1 = r_283_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_2_clock = clock;
  assign mesh_11_2_io_in_a_0 = r_178_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_2_io_in_a_1 = r_178_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_2_io_in_b_0 = pipe_b_43_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_b_1 = pipe_b_43_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_d_0 = pipe_b_299_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_d_1 = pipe_b_299_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_control_0_dataflow = mesh_11_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_control_0_propagate = mesh_11_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_control_0_shift = mesh_11_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_control_1_dataflow = mesh_11_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_control_1_propagate = mesh_11_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_control_1_shift = mesh_11_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_2_io_in_id_0 = r_555_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_2_io_in_id_1 = r_555_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_2_io_in_last_0 = r_811_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_2_io_in_last_1 = r_811_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_2_io_in_valid_0 = r_299_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_2_io_in_valid_1 = r_299_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_3_clock = clock;
  assign mesh_11_3_io_in_a_0 = r_179_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_3_io_in_a_1 = r_179_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_3_io_in_b_0 = pipe_b_59_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_b_1 = pipe_b_59_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_d_0 = pipe_b_315_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_d_1 = pipe_b_315_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_control_0_dataflow = mesh_11_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_control_0_propagate = mesh_11_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_control_0_shift = mesh_11_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_control_1_dataflow = mesh_11_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_control_1_propagate = mesh_11_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_control_1_shift = mesh_11_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_3_io_in_id_0 = r_571_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_3_io_in_id_1 = r_571_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_3_io_in_last_0 = r_827_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_3_io_in_last_1 = r_827_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_3_io_in_valid_0 = r_315_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_3_io_in_valid_1 = r_315_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_4_clock = clock;
  assign mesh_11_4_io_in_a_0 = r_180_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_4_io_in_a_1 = r_180_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_4_io_in_b_0 = pipe_b_75_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_b_1 = pipe_b_75_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_d_0 = pipe_b_331_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_d_1 = pipe_b_331_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_control_0_dataflow = mesh_11_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_control_0_propagate = mesh_11_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_control_0_shift = mesh_11_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_control_1_dataflow = mesh_11_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_control_1_propagate = mesh_11_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_control_1_shift = mesh_11_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_4_io_in_id_0 = r_587_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_4_io_in_id_1 = r_587_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_4_io_in_last_0 = r_843_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_4_io_in_last_1 = r_843_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_4_io_in_valid_0 = r_331_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_4_io_in_valid_1 = r_331_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_5_clock = clock;
  assign mesh_11_5_io_in_a_0 = r_181_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_5_io_in_a_1 = r_181_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_5_io_in_b_0 = pipe_b_91_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_b_1 = pipe_b_91_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_d_0 = pipe_b_347_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_d_1 = pipe_b_347_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_control_0_dataflow = mesh_11_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_control_0_propagate = mesh_11_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_control_0_shift = mesh_11_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_control_1_dataflow = mesh_11_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_control_1_propagate = mesh_11_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_control_1_shift = mesh_11_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_5_io_in_id_0 = r_603_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_5_io_in_id_1 = r_603_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_5_io_in_last_0 = r_859_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_5_io_in_last_1 = r_859_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_5_io_in_valid_0 = r_347_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_5_io_in_valid_1 = r_347_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_6_clock = clock;
  assign mesh_11_6_io_in_a_0 = r_182_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_6_io_in_a_1 = r_182_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_6_io_in_b_0 = pipe_b_107_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_b_1 = pipe_b_107_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_d_0 = pipe_b_363_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_d_1 = pipe_b_363_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_control_0_dataflow = mesh_11_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_control_0_propagate = mesh_11_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_control_0_shift = mesh_11_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_control_1_dataflow = mesh_11_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_control_1_propagate = mesh_11_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_control_1_shift = mesh_11_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_6_io_in_id_0 = r_619_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_6_io_in_id_1 = r_619_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_6_io_in_last_0 = r_875_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_6_io_in_last_1 = r_875_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_6_io_in_valid_0 = r_363_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_6_io_in_valid_1 = r_363_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_7_clock = clock;
  assign mesh_11_7_io_in_a_0 = r_183_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_7_io_in_a_1 = r_183_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_7_io_in_b_0 = pipe_b_123_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_b_1 = pipe_b_123_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_d_0 = pipe_b_379_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_d_1 = pipe_b_379_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_control_0_dataflow = mesh_11_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_control_0_propagate = mesh_11_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_control_0_shift = mesh_11_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_control_1_dataflow = mesh_11_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_control_1_propagate = mesh_11_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_control_1_shift = mesh_11_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_7_io_in_id_0 = r_635_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_7_io_in_id_1 = r_635_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_7_io_in_last_0 = r_891_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_7_io_in_last_1 = r_891_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_7_io_in_valid_0 = r_379_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_7_io_in_valid_1 = r_379_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_8_clock = clock;
  assign mesh_11_8_io_in_a_0 = r_184_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_8_io_in_a_1 = r_184_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_8_io_in_b_0 = pipe_b_139_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_b_1 = pipe_b_139_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_d_0 = pipe_b_395_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_d_1 = pipe_b_395_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_control_0_dataflow = mesh_11_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_control_0_propagate = mesh_11_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_control_0_shift = mesh_11_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_control_1_dataflow = mesh_11_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_control_1_propagate = mesh_11_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_control_1_shift = mesh_11_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_8_io_in_id_0 = r_651_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_8_io_in_id_1 = r_651_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_8_io_in_last_0 = r_907_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_8_io_in_last_1 = r_907_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_8_io_in_valid_0 = r_395_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_8_io_in_valid_1 = r_395_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_9_clock = clock;
  assign mesh_11_9_io_in_a_0 = r_185_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_9_io_in_a_1 = r_185_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_9_io_in_b_0 = pipe_b_155_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_b_1 = pipe_b_155_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_d_0 = pipe_b_411_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_d_1 = pipe_b_411_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_control_0_dataflow = mesh_11_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_control_0_propagate = mesh_11_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_control_0_shift = mesh_11_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_control_1_dataflow = mesh_11_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_control_1_propagate = mesh_11_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_control_1_shift = mesh_11_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_9_io_in_id_0 = r_667_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_9_io_in_id_1 = r_667_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_9_io_in_last_0 = r_923_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_9_io_in_last_1 = r_923_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_9_io_in_valid_0 = r_411_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_9_io_in_valid_1 = r_411_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_10_clock = clock;
  assign mesh_11_10_io_in_a_0 = r_186_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_10_io_in_a_1 = r_186_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_10_io_in_b_0 = pipe_b_171_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_b_1 = pipe_b_171_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_d_0 = pipe_b_427_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_d_1 = pipe_b_427_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_control_0_dataflow = mesh_11_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_control_0_propagate = mesh_11_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_control_0_shift = mesh_11_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_control_1_dataflow = mesh_11_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_control_1_propagate = mesh_11_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_control_1_shift = mesh_11_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_10_io_in_id_0 = r_683_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_10_io_in_id_1 = r_683_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_10_io_in_last_0 = r_939_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_10_io_in_last_1 = r_939_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_10_io_in_valid_0 = r_427_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_10_io_in_valid_1 = r_427_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_11_clock = clock;
  assign mesh_11_11_io_in_a_0 = r_187_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_11_io_in_a_1 = r_187_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_11_io_in_b_0 = pipe_b_187_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_b_1 = pipe_b_187_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_d_0 = pipe_b_443_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_d_1 = pipe_b_443_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_control_0_dataflow = mesh_11_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_control_0_propagate = mesh_11_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_control_0_shift = mesh_11_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_control_1_dataflow = mesh_11_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_control_1_propagate = mesh_11_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_control_1_shift = mesh_11_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_11_io_in_id_0 = r_699_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_11_io_in_id_1 = r_699_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_11_io_in_last_0 = r_955_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_11_io_in_last_1 = r_955_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_11_io_in_valid_0 = r_443_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_11_io_in_valid_1 = r_443_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_12_clock = clock;
  assign mesh_11_12_io_in_a_0 = r_188_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_12_io_in_a_1 = r_188_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_12_io_in_b_0 = pipe_b_203_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_b_1 = pipe_b_203_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_d_0 = pipe_b_459_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_d_1 = pipe_b_459_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_control_0_dataflow = mesh_11_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_control_0_propagate = mesh_11_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_control_0_shift = mesh_11_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_control_1_dataflow = mesh_11_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_control_1_propagate = mesh_11_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_control_1_shift = mesh_11_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_12_io_in_id_0 = r_715_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_12_io_in_id_1 = r_715_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_12_io_in_last_0 = r_971_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_12_io_in_last_1 = r_971_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_12_io_in_valid_0 = r_459_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_12_io_in_valid_1 = r_459_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_13_clock = clock;
  assign mesh_11_13_io_in_a_0 = r_189_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_13_io_in_a_1 = r_189_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_13_io_in_b_0 = pipe_b_219_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_b_1 = pipe_b_219_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_d_0 = pipe_b_475_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_d_1 = pipe_b_475_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_control_0_dataflow = mesh_11_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_control_0_propagate = mesh_11_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_control_0_shift = mesh_11_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_control_1_dataflow = mesh_11_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_control_1_propagate = mesh_11_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_control_1_shift = mesh_11_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_13_io_in_id_0 = r_731_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_13_io_in_id_1 = r_731_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_13_io_in_last_0 = r_987_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_13_io_in_last_1 = r_987_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_13_io_in_valid_0 = r_475_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_13_io_in_valid_1 = r_475_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_14_clock = clock;
  assign mesh_11_14_io_in_a_0 = r_190_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_14_io_in_a_1 = r_190_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_14_io_in_b_0 = pipe_b_235_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_b_1 = pipe_b_235_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_d_0 = pipe_b_491_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_d_1 = pipe_b_491_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_control_0_dataflow = mesh_11_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_control_0_propagate = mesh_11_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_control_0_shift = mesh_11_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_control_1_dataflow = mesh_11_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_control_1_propagate = mesh_11_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_control_1_shift = mesh_11_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_14_io_in_id_0 = r_747_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_14_io_in_id_1 = r_747_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_14_io_in_last_0 = r_1003_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_14_io_in_last_1 = r_1003_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_14_io_in_valid_0 = r_491_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_14_io_in_valid_1 = r_491_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_15_clock = clock;
  assign mesh_11_15_io_in_a_0 = r_191_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_15_io_in_a_1 = r_191_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_11_15_io_in_b_0 = pipe_b_251_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_b_1 = pipe_b_251_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_d_0 = pipe_b_507_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_d_1 = pipe_b_507_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_control_0_dataflow = mesh_11_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_control_0_propagate = mesh_11_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_control_0_shift = mesh_11_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_control_1_dataflow = mesh_11_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_control_1_propagate = mesh_11_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_control_1_shift = mesh_11_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_11_15_io_in_id_0 = r_763_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_15_io_in_id_1 = r_763_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_11_15_io_in_last_0 = r_1019_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_15_io_in_last_1 = r_1019_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_11_15_io_in_valid_0 = r_507_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_11_15_io_in_valid_1 = r_507_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_0_clock = clock;
  assign mesh_12_0_io_in_a_0 = r_192_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_0_io_in_a_1 = r_192_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_0_io_in_b_0 = pipe_b_12_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_b_1 = pipe_b_12_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_d_0 = pipe_b_268_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_d_1 = pipe_b_268_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_control_0_dataflow = mesh_12_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_control_0_propagate = mesh_12_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_control_0_shift = mesh_12_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_control_1_dataflow = mesh_12_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_control_1_propagate = mesh_12_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_control_1_shift = mesh_12_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_0_io_in_id_0 = r_524_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_0_io_in_id_1 = r_524_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_0_io_in_last_0 = r_780_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_0_io_in_last_1 = r_780_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_0_io_in_valid_0 = r_268_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_0_io_in_valid_1 = r_268_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_1_clock = clock;
  assign mesh_12_1_io_in_a_0 = r_193_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_1_io_in_a_1 = r_193_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_1_io_in_b_0 = pipe_b_28_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_b_1 = pipe_b_28_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_d_0 = pipe_b_284_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_d_1 = pipe_b_284_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_control_0_dataflow = mesh_12_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_control_0_propagate = mesh_12_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_control_0_shift = mesh_12_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_control_1_dataflow = mesh_12_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_control_1_propagate = mesh_12_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_control_1_shift = mesh_12_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_1_io_in_id_0 = r_540_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_1_io_in_id_1 = r_540_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_1_io_in_last_0 = r_796_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_1_io_in_last_1 = r_796_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_1_io_in_valid_0 = r_284_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_1_io_in_valid_1 = r_284_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_2_clock = clock;
  assign mesh_12_2_io_in_a_0 = r_194_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_2_io_in_a_1 = r_194_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_2_io_in_b_0 = pipe_b_44_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_b_1 = pipe_b_44_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_d_0 = pipe_b_300_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_d_1 = pipe_b_300_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_control_0_dataflow = mesh_12_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_control_0_propagate = mesh_12_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_control_0_shift = mesh_12_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_control_1_dataflow = mesh_12_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_control_1_propagate = mesh_12_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_control_1_shift = mesh_12_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_2_io_in_id_0 = r_556_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_2_io_in_id_1 = r_556_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_2_io_in_last_0 = r_812_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_2_io_in_last_1 = r_812_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_2_io_in_valid_0 = r_300_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_2_io_in_valid_1 = r_300_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_3_clock = clock;
  assign mesh_12_3_io_in_a_0 = r_195_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_3_io_in_a_1 = r_195_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_3_io_in_b_0 = pipe_b_60_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_b_1 = pipe_b_60_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_d_0 = pipe_b_316_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_d_1 = pipe_b_316_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_control_0_dataflow = mesh_12_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_control_0_propagate = mesh_12_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_control_0_shift = mesh_12_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_control_1_dataflow = mesh_12_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_control_1_propagate = mesh_12_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_control_1_shift = mesh_12_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_3_io_in_id_0 = r_572_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_3_io_in_id_1 = r_572_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_3_io_in_last_0 = r_828_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_3_io_in_last_1 = r_828_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_3_io_in_valid_0 = r_316_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_3_io_in_valid_1 = r_316_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_4_clock = clock;
  assign mesh_12_4_io_in_a_0 = r_196_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_4_io_in_a_1 = r_196_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_4_io_in_b_0 = pipe_b_76_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_b_1 = pipe_b_76_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_d_0 = pipe_b_332_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_d_1 = pipe_b_332_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_control_0_dataflow = mesh_12_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_control_0_propagate = mesh_12_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_control_0_shift = mesh_12_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_control_1_dataflow = mesh_12_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_control_1_propagate = mesh_12_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_control_1_shift = mesh_12_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_4_io_in_id_0 = r_588_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_4_io_in_id_1 = r_588_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_4_io_in_last_0 = r_844_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_4_io_in_last_1 = r_844_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_4_io_in_valid_0 = r_332_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_4_io_in_valid_1 = r_332_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_5_clock = clock;
  assign mesh_12_5_io_in_a_0 = r_197_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_5_io_in_a_1 = r_197_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_5_io_in_b_0 = pipe_b_92_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_b_1 = pipe_b_92_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_d_0 = pipe_b_348_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_d_1 = pipe_b_348_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_control_0_dataflow = mesh_12_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_control_0_propagate = mesh_12_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_control_0_shift = mesh_12_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_control_1_dataflow = mesh_12_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_control_1_propagate = mesh_12_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_control_1_shift = mesh_12_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_5_io_in_id_0 = r_604_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_5_io_in_id_1 = r_604_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_5_io_in_last_0 = r_860_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_5_io_in_last_1 = r_860_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_5_io_in_valid_0 = r_348_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_5_io_in_valid_1 = r_348_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_6_clock = clock;
  assign mesh_12_6_io_in_a_0 = r_198_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_6_io_in_a_1 = r_198_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_6_io_in_b_0 = pipe_b_108_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_b_1 = pipe_b_108_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_d_0 = pipe_b_364_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_d_1 = pipe_b_364_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_control_0_dataflow = mesh_12_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_control_0_propagate = mesh_12_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_control_0_shift = mesh_12_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_control_1_dataflow = mesh_12_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_control_1_propagate = mesh_12_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_control_1_shift = mesh_12_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_6_io_in_id_0 = r_620_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_6_io_in_id_1 = r_620_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_6_io_in_last_0 = r_876_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_6_io_in_last_1 = r_876_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_6_io_in_valid_0 = r_364_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_6_io_in_valid_1 = r_364_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_7_clock = clock;
  assign mesh_12_7_io_in_a_0 = r_199_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_7_io_in_a_1 = r_199_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_7_io_in_b_0 = pipe_b_124_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_b_1 = pipe_b_124_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_d_0 = pipe_b_380_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_d_1 = pipe_b_380_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_control_0_dataflow = mesh_12_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_control_0_propagate = mesh_12_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_control_0_shift = mesh_12_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_control_1_dataflow = mesh_12_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_control_1_propagate = mesh_12_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_control_1_shift = mesh_12_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_7_io_in_id_0 = r_636_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_7_io_in_id_1 = r_636_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_7_io_in_last_0 = r_892_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_7_io_in_last_1 = r_892_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_7_io_in_valid_0 = r_380_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_7_io_in_valid_1 = r_380_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_8_clock = clock;
  assign mesh_12_8_io_in_a_0 = r_200_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_8_io_in_a_1 = r_200_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_8_io_in_b_0 = pipe_b_140_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_b_1 = pipe_b_140_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_d_0 = pipe_b_396_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_d_1 = pipe_b_396_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_control_0_dataflow = mesh_12_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_control_0_propagate = mesh_12_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_control_0_shift = mesh_12_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_control_1_dataflow = mesh_12_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_control_1_propagate = mesh_12_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_control_1_shift = mesh_12_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_8_io_in_id_0 = r_652_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_8_io_in_id_1 = r_652_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_8_io_in_last_0 = r_908_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_8_io_in_last_1 = r_908_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_8_io_in_valid_0 = r_396_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_8_io_in_valid_1 = r_396_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_9_clock = clock;
  assign mesh_12_9_io_in_a_0 = r_201_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_9_io_in_a_1 = r_201_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_9_io_in_b_0 = pipe_b_156_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_b_1 = pipe_b_156_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_d_0 = pipe_b_412_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_d_1 = pipe_b_412_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_control_0_dataflow = mesh_12_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_control_0_propagate = mesh_12_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_control_0_shift = mesh_12_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_control_1_dataflow = mesh_12_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_control_1_propagate = mesh_12_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_control_1_shift = mesh_12_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_9_io_in_id_0 = r_668_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_9_io_in_id_1 = r_668_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_9_io_in_last_0 = r_924_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_9_io_in_last_1 = r_924_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_9_io_in_valid_0 = r_412_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_9_io_in_valid_1 = r_412_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_10_clock = clock;
  assign mesh_12_10_io_in_a_0 = r_202_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_10_io_in_a_1 = r_202_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_10_io_in_b_0 = pipe_b_172_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_b_1 = pipe_b_172_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_d_0 = pipe_b_428_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_d_1 = pipe_b_428_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_control_0_dataflow = mesh_12_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_control_0_propagate = mesh_12_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_control_0_shift = mesh_12_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_control_1_dataflow = mesh_12_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_control_1_propagate = mesh_12_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_control_1_shift = mesh_12_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_10_io_in_id_0 = r_684_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_10_io_in_id_1 = r_684_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_10_io_in_last_0 = r_940_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_10_io_in_last_1 = r_940_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_10_io_in_valid_0 = r_428_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_10_io_in_valid_1 = r_428_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_11_clock = clock;
  assign mesh_12_11_io_in_a_0 = r_203_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_11_io_in_a_1 = r_203_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_11_io_in_b_0 = pipe_b_188_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_b_1 = pipe_b_188_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_d_0 = pipe_b_444_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_d_1 = pipe_b_444_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_control_0_dataflow = mesh_12_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_control_0_propagate = mesh_12_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_control_0_shift = mesh_12_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_control_1_dataflow = mesh_12_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_control_1_propagate = mesh_12_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_control_1_shift = mesh_12_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_11_io_in_id_0 = r_700_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_11_io_in_id_1 = r_700_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_11_io_in_last_0 = r_956_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_11_io_in_last_1 = r_956_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_11_io_in_valid_0 = r_444_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_11_io_in_valid_1 = r_444_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_12_clock = clock;
  assign mesh_12_12_io_in_a_0 = r_204_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_12_io_in_a_1 = r_204_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_12_io_in_b_0 = pipe_b_204_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_b_1 = pipe_b_204_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_d_0 = pipe_b_460_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_d_1 = pipe_b_460_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_control_0_dataflow = mesh_12_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_control_0_propagate = mesh_12_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_control_0_shift = mesh_12_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_control_1_dataflow = mesh_12_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_control_1_propagate = mesh_12_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_control_1_shift = mesh_12_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_12_io_in_id_0 = r_716_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_12_io_in_id_1 = r_716_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_12_io_in_last_0 = r_972_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_12_io_in_last_1 = r_972_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_12_io_in_valid_0 = r_460_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_12_io_in_valid_1 = r_460_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_13_clock = clock;
  assign mesh_12_13_io_in_a_0 = r_205_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_13_io_in_a_1 = r_205_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_13_io_in_b_0 = pipe_b_220_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_b_1 = pipe_b_220_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_d_0 = pipe_b_476_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_d_1 = pipe_b_476_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_control_0_dataflow = mesh_12_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_control_0_propagate = mesh_12_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_control_0_shift = mesh_12_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_control_1_dataflow = mesh_12_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_control_1_propagate = mesh_12_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_control_1_shift = mesh_12_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_13_io_in_id_0 = r_732_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_13_io_in_id_1 = r_732_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_13_io_in_last_0 = r_988_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_13_io_in_last_1 = r_988_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_13_io_in_valid_0 = r_476_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_13_io_in_valid_1 = r_476_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_14_clock = clock;
  assign mesh_12_14_io_in_a_0 = r_206_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_14_io_in_a_1 = r_206_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_14_io_in_b_0 = pipe_b_236_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_b_1 = pipe_b_236_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_d_0 = pipe_b_492_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_d_1 = pipe_b_492_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_control_0_dataflow = mesh_12_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_control_0_propagate = mesh_12_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_control_0_shift = mesh_12_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_control_1_dataflow = mesh_12_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_control_1_propagate = mesh_12_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_control_1_shift = mesh_12_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_14_io_in_id_0 = r_748_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_14_io_in_id_1 = r_748_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_14_io_in_last_0 = r_1004_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_14_io_in_last_1 = r_1004_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_14_io_in_valid_0 = r_492_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_14_io_in_valid_1 = r_492_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_15_clock = clock;
  assign mesh_12_15_io_in_a_0 = r_207_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_15_io_in_a_1 = r_207_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_12_15_io_in_b_0 = pipe_b_252_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_b_1 = pipe_b_252_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_d_0 = pipe_b_508_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_d_1 = pipe_b_508_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_control_0_dataflow = mesh_12_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_control_0_propagate = mesh_12_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_control_0_shift = mesh_12_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_control_1_dataflow = mesh_12_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_control_1_propagate = mesh_12_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_control_1_shift = mesh_12_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_12_15_io_in_id_0 = r_764_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_15_io_in_id_1 = r_764_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_12_15_io_in_last_0 = r_1020_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_15_io_in_last_1 = r_1020_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_12_15_io_in_valid_0 = r_508_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_12_15_io_in_valid_1 = r_508_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_0_clock = clock;
  assign mesh_13_0_io_in_a_0 = r_208_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_0_io_in_a_1 = r_208_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_0_io_in_b_0 = pipe_b_13_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_b_1 = pipe_b_13_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_d_0 = pipe_b_269_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_d_1 = pipe_b_269_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_control_0_dataflow = mesh_13_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_control_0_propagate = mesh_13_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_control_0_shift = mesh_13_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_control_1_dataflow = mesh_13_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_control_1_propagate = mesh_13_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_control_1_shift = mesh_13_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_0_io_in_id_0 = r_525_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_0_io_in_id_1 = r_525_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_0_io_in_last_0 = r_781_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_0_io_in_last_1 = r_781_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_0_io_in_valid_0 = r_269_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_0_io_in_valid_1 = r_269_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_1_clock = clock;
  assign mesh_13_1_io_in_a_0 = r_209_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_1_io_in_a_1 = r_209_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_1_io_in_b_0 = pipe_b_29_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_b_1 = pipe_b_29_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_d_0 = pipe_b_285_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_d_1 = pipe_b_285_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_control_0_dataflow = mesh_13_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_control_0_propagate = mesh_13_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_control_0_shift = mesh_13_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_control_1_dataflow = mesh_13_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_control_1_propagate = mesh_13_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_control_1_shift = mesh_13_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_1_io_in_id_0 = r_541_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_1_io_in_id_1 = r_541_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_1_io_in_last_0 = r_797_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_1_io_in_last_1 = r_797_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_1_io_in_valid_0 = r_285_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_1_io_in_valid_1 = r_285_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_2_clock = clock;
  assign mesh_13_2_io_in_a_0 = r_210_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_2_io_in_a_1 = r_210_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_2_io_in_b_0 = pipe_b_45_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_b_1 = pipe_b_45_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_d_0 = pipe_b_301_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_d_1 = pipe_b_301_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_control_0_dataflow = mesh_13_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_control_0_propagate = mesh_13_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_control_0_shift = mesh_13_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_control_1_dataflow = mesh_13_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_control_1_propagate = mesh_13_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_control_1_shift = mesh_13_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_2_io_in_id_0 = r_557_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_2_io_in_id_1 = r_557_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_2_io_in_last_0 = r_813_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_2_io_in_last_1 = r_813_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_2_io_in_valid_0 = r_301_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_2_io_in_valid_1 = r_301_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_3_clock = clock;
  assign mesh_13_3_io_in_a_0 = r_211_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_3_io_in_a_1 = r_211_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_3_io_in_b_0 = pipe_b_61_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_b_1 = pipe_b_61_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_d_0 = pipe_b_317_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_d_1 = pipe_b_317_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_control_0_dataflow = mesh_13_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_control_0_propagate = mesh_13_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_control_0_shift = mesh_13_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_control_1_dataflow = mesh_13_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_control_1_propagate = mesh_13_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_control_1_shift = mesh_13_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_3_io_in_id_0 = r_573_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_3_io_in_id_1 = r_573_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_3_io_in_last_0 = r_829_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_3_io_in_last_1 = r_829_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_3_io_in_valid_0 = r_317_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_3_io_in_valid_1 = r_317_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_4_clock = clock;
  assign mesh_13_4_io_in_a_0 = r_212_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_4_io_in_a_1 = r_212_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_4_io_in_b_0 = pipe_b_77_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_b_1 = pipe_b_77_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_d_0 = pipe_b_333_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_d_1 = pipe_b_333_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_control_0_dataflow = mesh_13_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_control_0_propagate = mesh_13_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_control_0_shift = mesh_13_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_control_1_dataflow = mesh_13_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_control_1_propagate = mesh_13_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_control_1_shift = mesh_13_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_4_io_in_id_0 = r_589_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_4_io_in_id_1 = r_589_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_4_io_in_last_0 = r_845_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_4_io_in_last_1 = r_845_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_4_io_in_valid_0 = r_333_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_4_io_in_valid_1 = r_333_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_5_clock = clock;
  assign mesh_13_5_io_in_a_0 = r_213_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_5_io_in_a_1 = r_213_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_5_io_in_b_0 = pipe_b_93_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_b_1 = pipe_b_93_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_d_0 = pipe_b_349_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_d_1 = pipe_b_349_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_control_0_dataflow = mesh_13_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_control_0_propagate = mesh_13_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_control_0_shift = mesh_13_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_control_1_dataflow = mesh_13_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_control_1_propagate = mesh_13_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_control_1_shift = mesh_13_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_5_io_in_id_0 = r_605_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_5_io_in_id_1 = r_605_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_5_io_in_last_0 = r_861_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_5_io_in_last_1 = r_861_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_5_io_in_valid_0 = r_349_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_5_io_in_valid_1 = r_349_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_6_clock = clock;
  assign mesh_13_6_io_in_a_0 = r_214_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_6_io_in_a_1 = r_214_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_6_io_in_b_0 = pipe_b_109_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_b_1 = pipe_b_109_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_d_0 = pipe_b_365_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_d_1 = pipe_b_365_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_control_0_dataflow = mesh_13_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_control_0_propagate = mesh_13_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_control_0_shift = mesh_13_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_control_1_dataflow = mesh_13_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_control_1_propagate = mesh_13_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_control_1_shift = mesh_13_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_6_io_in_id_0 = r_621_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_6_io_in_id_1 = r_621_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_6_io_in_last_0 = r_877_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_6_io_in_last_1 = r_877_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_6_io_in_valid_0 = r_365_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_6_io_in_valid_1 = r_365_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_7_clock = clock;
  assign mesh_13_7_io_in_a_0 = r_215_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_7_io_in_a_1 = r_215_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_7_io_in_b_0 = pipe_b_125_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_b_1 = pipe_b_125_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_d_0 = pipe_b_381_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_d_1 = pipe_b_381_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_control_0_dataflow = mesh_13_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_control_0_propagate = mesh_13_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_control_0_shift = mesh_13_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_control_1_dataflow = mesh_13_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_control_1_propagate = mesh_13_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_control_1_shift = mesh_13_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_7_io_in_id_0 = r_637_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_7_io_in_id_1 = r_637_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_7_io_in_last_0 = r_893_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_7_io_in_last_1 = r_893_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_7_io_in_valid_0 = r_381_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_7_io_in_valid_1 = r_381_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_8_clock = clock;
  assign mesh_13_8_io_in_a_0 = r_216_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_8_io_in_a_1 = r_216_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_8_io_in_b_0 = pipe_b_141_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_b_1 = pipe_b_141_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_d_0 = pipe_b_397_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_d_1 = pipe_b_397_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_control_0_dataflow = mesh_13_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_control_0_propagate = mesh_13_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_control_0_shift = mesh_13_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_control_1_dataflow = mesh_13_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_control_1_propagate = mesh_13_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_control_1_shift = mesh_13_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_8_io_in_id_0 = r_653_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_8_io_in_id_1 = r_653_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_8_io_in_last_0 = r_909_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_8_io_in_last_1 = r_909_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_8_io_in_valid_0 = r_397_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_8_io_in_valid_1 = r_397_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_9_clock = clock;
  assign mesh_13_9_io_in_a_0 = r_217_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_9_io_in_a_1 = r_217_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_9_io_in_b_0 = pipe_b_157_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_b_1 = pipe_b_157_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_d_0 = pipe_b_413_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_d_1 = pipe_b_413_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_control_0_dataflow = mesh_13_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_control_0_propagate = mesh_13_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_control_0_shift = mesh_13_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_control_1_dataflow = mesh_13_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_control_1_propagate = mesh_13_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_control_1_shift = mesh_13_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_9_io_in_id_0 = r_669_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_9_io_in_id_1 = r_669_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_9_io_in_last_0 = r_925_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_9_io_in_last_1 = r_925_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_9_io_in_valid_0 = r_413_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_9_io_in_valid_1 = r_413_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_10_clock = clock;
  assign mesh_13_10_io_in_a_0 = r_218_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_10_io_in_a_1 = r_218_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_10_io_in_b_0 = pipe_b_173_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_b_1 = pipe_b_173_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_d_0 = pipe_b_429_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_d_1 = pipe_b_429_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_control_0_dataflow = mesh_13_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_control_0_propagate = mesh_13_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_control_0_shift = mesh_13_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_control_1_dataflow = mesh_13_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_control_1_propagate = mesh_13_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_control_1_shift = mesh_13_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_10_io_in_id_0 = r_685_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_10_io_in_id_1 = r_685_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_10_io_in_last_0 = r_941_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_10_io_in_last_1 = r_941_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_10_io_in_valid_0 = r_429_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_10_io_in_valid_1 = r_429_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_11_clock = clock;
  assign mesh_13_11_io_in_a_0 = r_219_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_11_io_in_a_1 = r_219_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_11_io_in_b_0 = pipe_b_189_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_b_1 = pipe_b_189_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_d_0 = pipe_b_445_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_d_1 = pipe_b_445_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_control_0_dataflow = mesh_13_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_control_0_propagate = mesh_13_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_control_0_shift = mesh_13_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_control_1_dataflow = mesh_13_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_control_1_propagate = mesh_13_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_control_1_shift = mesh_13_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_11_io_in_id_0 = r_701_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_11_io_in_id_1 = r_701_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_11_io_in_last_0 = r_957_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_11_io_in_last_1 = r_957_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_11_io_in_valid_0 = r_445_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_11_io_in_valid_1 = r_445_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_12_clock = clock;
  assign mesh_13_12_io_in_a_0 = r_220_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_12_io_in_a_1 = r_220_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_12_io_in_b_0 = pipe_b_205_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_b_1 = pipe_b_205_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_d_0 = pipe_b_461_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_d_1 = pipe_b_461_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_control_0_dataflow = mesh_13_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_control_0_propagate = mesh_13_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_control_0_shift = mesh_13_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_control_1_dataflow = mesh_13_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_control_1_propagate = mesh_13_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_control_1_shift = mesh_13_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_12_io_in_id_0 = r_717_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_12_io_in_id_1 = r_717_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_12_io_in_last_0 = r_973_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_12_io_in_last_1 = r_973_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_12_io_in_valid_0 = r_461_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_12_io_in_valid_1 = r_461_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_13_clock = clock;
  assign mesh_13_13_io_in_a_0 = r_221_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_13_io_in_a_1 = r_221_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_13_io_in_b_0 = pipe_b_221_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_b_1 = pipe_b_221_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_d_0 = pipe_b_477_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_d_1 = pipe_b_477_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_control_0_dataflow = mesh_13_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_control_0_propagate = mesh_13_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_control_0_shift = mesh_13_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_control_1_dataflow = mesh_13_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_control_1_propagate = mesh_13_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_control_1_shift = mesh_13_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_13_io_in_id_0 = r_733_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_13_io_in_id_1 = r_733_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_13_io_in_last_0 = r_989_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_13_io_in_last_1 = r_989_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_13_io_in_valid_0 = r_477_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_13_io_in_valid_1 = r_477_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_14_clock = clock;
  assign mesh_13_14_io_in_a_0 = r_222_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_14_io_in_a_1 = r_222_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_14_io_in_b_0 = pipe_b_237_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_b_1 = pipe_b_237_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_d_0 = pipe_b_493_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_d_1 = pipe_b_493_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_control_0_dataflow = mesh_13_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_control_0_propagate = mesh_13_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_control_0_shift = mesh_13_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_control_1_dataflow = mesh_13_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_control_1_propagate = mesh_13_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_control_1_shift = mesh_13_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_14_io_in_id_0 = r_749_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_14_io_in_id_1 = r_749_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_14_io_in_last_0 = r_1005_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_14_io_in_last_1 = r_1005_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_14_io_in_valid_0 = r_493_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_14_io_in_valid_1 = r_493_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_15_clock = clock;
  assign mesh_13_15_io_in_a_0 = r_223_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_15_io_in_a_1 = r_223_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_13_15_io_in_b_0 = pipe_b_253_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_b_1 = pipe_b_253_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_d_0 = pipe_b_509_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_d_1 = pipe_b_509_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_control_0_dataflow = mesh_13_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_control_0_propagate = mesh_13_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_control_0_shift = mesh_13_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_control_1_dataflow = mesh_13_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_control_1_propagate = mesh_13_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_control_1_shift = mesh_13_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_13_15_io_in_id_0 = r_765_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_15_io_in_id_1 = r_765_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_13_15_io_in_last_0 = r_1021_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_15_io_in_last_1 = r_1021_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_13_15_io_in_valid_0 = r_509_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_13_15_io_in_valid_1 = r_509_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_0_clock = clock;
  assign mesh_14_0_io_in_a_0 = r_224_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_0_io_in_a_1 = r_224_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_0_io_in_b_0 = pipe_b_14_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_b_1 = pipe_b_14_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_d_0 = pipe_b_270_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_d_1 = pipe_b_270_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_control_0_dataflow = mesh_14_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_control_0_propagate = mesh_14_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_control_0_shift = mesh_14_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_control_1_dataflow = mesh_14_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_control_1_propagate = mesh_14_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_control_1_shift = mesh_14_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_0_io_in_id_0 = r_526_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_0_io_in_id_1 = r_526_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_0_io_in_last_0 = r_782_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_0_io_in_last_1 = r_782_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_0_io_in_valid_0 = r_270_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_0_io_in_valid_1 = r_270_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_1_clock = clock;
  assign mesh_14_1_io_in_a_0 = r_225_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_1_io_in_a_1 = r_225_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_1_io_in_b_0 = pipe_b_30_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_b_1 = pipe_b_30_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_d_0 = pipe_b_286_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_d_1 = pipe_b_286_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_control_0_dataflow = mesh_14_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_control_0_propagate = mesh_14_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_control_0_shift = mesh_14_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_control_1_dataflow = mesh_14_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_control_1_propagate = mesh_14_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_control_1_shift = mesh_14_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_1_io_in_id_0 = r_542_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_1_io_in_id_1 = r_542_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_1_io_in_last_0 = r_798_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_1_io_in_last_1 = r_798_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_1_io_in_valid_0 = r_286_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_1_io_in_valid_1 = r_286_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_2_clock = clock;
  assign mesh_14_2_io_in_a_0 = r_226_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_2_io_in_a_1 = r_226_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_2_io_in_b_0 = pipe_b_46_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_b_1 = pipe_b_46_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_d_0 = pipe_b_302_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_d_1 = pipe_b_302_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_control_0_dataflow = mesh_14_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_control_0_propagate = mesh_14_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_control_0_shift = mesh_14_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_control_1_dataflow = mesh_14_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_control_1_propagate = mesh_14_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_control_1_shift = mesh_14_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_2_io_in_id_0 = r_558_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_2_io_in_id_1 = r_558_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_2_io_in_last_0 = r_814_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_2_io_in_last_1 = r_814_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_2_io_in_valid_0 = r_302_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_2_io_in_valid_1 = r_302_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_3_clock = clock;
  assign mesh_14_3_io_in_a_0 = r_227_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_3_io_in_a_1 = r_227_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_3_io_in_b_0 = pipe_b_62_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_b_1 = pipe_b_62_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_d_0 = pipe_b_318_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_d_1 = pipe_b_318_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_control_0_dataflow = mesh_14_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_control_0_propagate = mesh_14_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_control_0_shift = mesh_14_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_control_1_dataflow = mesh_14_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_control_1_propagate = mesh_14_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_control_1_shift = mesh_14_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_3_io_in_id_0 = r_574_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_3_io_in_id_1 = r_574_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_3_io_in_last_0 = r_830_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_3_io_in_last_1 = r_830_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_3_io_in_valid_0 = r_318_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_3_io_in_valid_1 = r_318_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_4_clock = clock;
  assign mesh_14_4_io_in_a_0 = r_228_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_4_io_in_a_1 = r_228_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_4_io_in_b_0 = pipe_b_78_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_b_1 = pipe_b_78_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_d_0 = pipe_b_334_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_d_1 = pipe_b_334_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_control_0_dataflow = mesh_14_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_control_0_propagate = mesh_14_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_control_0_shift = mesh_14_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_control_1_dataflow = mesh_14_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_control_1_propagate = mesh_14_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_control_1_shift = mesh_14_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_4_io_in_id_0 = r_590_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_4_io_in_id_1 = r_590_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_4_io_in_last_0 = r_846_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_4_io_in_last_1 = r_846_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_4_io_in_valid_0 = r_334_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_4_io_in_valid_1 = r_334_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_5_clock = clock;
  assign mesh_14_5_io_in_a_0 = r_229_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_5_io_in_a_1 = r_229_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_5_io_in_b_0 = pipe_b_94_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_b_1 = pipe_b_94_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_d_0 = pipe_b_350_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_d_1 = pipe_b_350_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_control_0_dataflow = mesh_14_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_control_0_propagate = mesh_14_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_control_0_shift = mesh_14_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_control_1_dataflow = mesh_14_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_control_1_propagate = mesh_14_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_control_1_shift = mesh_14_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_5_io_in_id_0 = r_606_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_5_io_in_id_1 = r_606_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_5_io_in_last_0 = r_862_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_5_io_in_last_1 = r_862_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_5_io_in_valid_0 = r_350_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_5_io_in_valid_1 = r_350_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_6_clock = clock;
  assign mesh_14_6_io_in_a_0 = r_230_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_6_io_in_a_1 = r_230_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_6_io_in_b_0 = pipe_b_110_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_b_1 = pipe_b_110_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_d_0 = pipe_b_366_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_d_1 = pipe_b_366_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_control_0_dataflow = mesh_14_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_control_0_propagate = mesh_14_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_control_0_shift = mesh_14_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_control_1_dataflow = mesh_14_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_control_1_propagate = mesh_14_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_control_1_shift = mesh_14_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_6_io_in_id_0 = r_622_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_6_io_in_id_1 = r_622_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_6_io_in_last_0 = r_878_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_6_io_in_last_1 = r_878_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_6_io_in_valid_0 = r_366_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_6_io_in_valid_1 = r_366_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_7_clock = clock;
  assign mesh_14_7_io_in_a_0 = r_231_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_7_io_in_a_1 = r_231_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_7_io_in_b_0 = pipe_b_126_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_b_1 = pipe_b_126_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_d_0 = pipe_b_382_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_d_1 = pipe_b_382_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_control_0_dataflow = mesh_14_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_control_0_propagate = mesh_14_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_control_0_shift = mesh_14_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_control_1_dataflow = mesh_14_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_control_1_propagate = mesh_14_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_control_1_shift = mesh_14_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_7_io_in_id_0 = r_638_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_7_io_in_id_1 = r_638_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_7_io_in_last_0 = r_894_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_7_io_in_last_1 = r_894_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_7_io_in_valid_0 = r_382_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_7_io_in_valid_1 = r_382_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_8_clock = clock;
  assign mesh_14_8_io_in_a_0 = r_232_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_8_io_in_a_1 = r_232_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_8_io_in_b_0 = pipe_b_142_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_b_1 = pipe_b_142_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_d_0 = pipe_b_398_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_d_1 = pipe_b_398_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_control_0_dataflow = mesh_14_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_control_0_propagate = mesh_14_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_control_0_shift = mesh_14_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_control_1_dataflow = mesh_14_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_control_1_propagate = mesh_14_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_control_1_shift = mesh_14_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_8_io_in_id_0 = r_654_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_8_io_in_id_1 = r_654_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_8_io_in_last_0 = r_910_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_8_io_in_last_1 = r_910_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_8_io_in_valid_0 = r_398_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_8_io_in_valid_1 = r_398_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_9_clock = clock;
  assign mesh_14_9_io_in_a_0 = r_233_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_9_io_in_a_1 = r_233_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_9_io_in_b_0 = pipe_b_158_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_b_1 = pipe_b_158_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_d_0 = pipe_b_414_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_d_1 = pipe_b_414_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_control_0_dataflow = mesh_14_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_control_0_propagate = mesh_14_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_control_0_shift = mesh_14_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_control_1_dataflow = mesh_14_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_control_1_propagate = mesh_14_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_control_1_shift = mesh_14_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_9_io_in_id_0 = r_670_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_9_io_in_id_1 = r_670_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_9_io_in_last_0 = r_926_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_9_io_in_last_1 = r_926_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_9_io_in_valid_0 = r_414_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_9_io_in_valid_1 = r_414_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_10_clock = clock;
  assign mesh_14_10_io_in_a_0 = r_234_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_10_io_in_a_1 = r_234_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_10_io_in_b_0 = pipe_b_174_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_b_1 = pipe_b_174_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_d_0 = pipe_b_430_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_d_1 = pipe_b_430_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_control_0_dataflow = mesh_14_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_control_0_propagate = mesh_14_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_control_0_shift = mesh_14_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_control_1_dataflow = mesh_14_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_control_1_propagate = mesh_14_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_control_1_shift = mesh_14_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_10_io_in_id_0 = r_686_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_10_io_in_id_1 = r_686_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_10_io_in_last_0 = r_942_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_10_io_in_last_1 = r_942_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_10_io_in_valid_0 = r_430_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_10_io_in_valid_1 = r_430_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_11_clock = clock;
  assign mesh_14_11_io_in_a_0 = r_235_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_11_io_in_a_1 = r_235_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_11_io_in_b_0 = pipe_b_190_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_b_1 = pipe_b_190_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_d_0 = pipe_b_446_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_d_1 = pipe_b_446_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_control_0_dataflow = mesh_14_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_control_0_propagate = mesh_14_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_control_0_shift = mesh_14_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_control_1_dataflow = mesh_14_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_control_1_propagate = mesh_14_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_control_1_shift = mesh_14_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_11_io_in_id_0 = r_702_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_11_io_in_id_1 = r_702_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_11_io_in_last_0 = r_958_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_11_io_in_last_1 = r_958_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_11_io_in_valid_0 = r_446_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_11_io_in_valid_1 = r_446_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_12_clock = clock;
  assign mesh_14_12_io_in_a_0 = r_236_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_12_io_in_a_1 = r_236_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_12_io_in_b_0 = pipe_b_206_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_b_1 = pipe_b_206_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_d_0 = pipe_b_462_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_d_1 = pipe_b_462_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_control_0_dataflow = mesh_14_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_control_0_propagate = mesh_14_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_control_0_shift = mesh_14_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_control_1_dataflow = mesh_14_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_control_1_propagate = mesh_14_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_control_1_shift = mesh_14_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_12_io_in_id_0 = r_718_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_12_io_in_id_1 = r_718_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_12_io_in_last_0 = r_974_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_12_io_in_last_1 = r_974_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_12_io_in_valid_0 = r_462_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_12_io_in_valid_1 = r_462_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_13_clock = clock;
  assign mesh_14_13_io_in_a_0 = r_237_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_13_io_in_a_1 = r_237_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_13_io_in_b_0 = pipe_b_222_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_b_1 = pipe_b_222_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_d_0 = pipe_b_478_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_d_1 = pipe_b_478_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_control_0_dataflow = mesh_14_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_control_0_propagate = mesh_14_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_control_0_shift = mesh_14_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_control_1_dataflow = mesh_14_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_control_1_propagate = mesh_14_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_control_1_shift = mesh_14_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_13_io_in_id_0 = r_734_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_13_io_in_id_1 = r_734_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_13_io_in_last_0 = r_990_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_13_io_in_last_1 = r_990_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_13_io_in_valid_0 = r_478_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_13_io_in_valid_1 = r_478_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_14_clock = clock;
  assign mesh_14_14_io_in_a_0 = r_238_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_14_io_in_a_1 = r_238_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_14_io_in_b_0 = pipe_b_238_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_b_1 = pipe_b_238_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_d_0 = pipe_b_494_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_d_1 = pipe_b_494_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_control_0_dataflow = mesh_14_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_control_0_propagate = mesh_14_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_control_0_shift = mesh_14_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_control_1_dataflow = mesh_14_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_control_1_propagate = mesh_14_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_control_1_shift = mesh_14_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_14_io_in_id_0 = r_750_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_14_io_in_id_1 = r_750_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_14_io_in_last_0 = r_1006_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_14_io_in_last_1 = r_1006_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_14_io_in_valid_0 = r_494_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_14_io_in_valid_1 = r_494_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_15_clock = clock;
  assign mesh_14_15_io_in_a_0 = r_239_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_15_io_in_a_1 = r_239_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_14_15_io_in_b_0 = pipe_b_254_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_b_1 = pipe_b_254_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_d_0 = pipe_b_510_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_d_1 = pipe_b_510_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_control_0_dataflow = mesh_14_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_control_0_propagate = mesh_14_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_control_0_shift = mesh_14_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_control_1_dataflow = mesh_14_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_control_1_propagate = mesh_14_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_control_1_shift = mesh_14_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_14_15_io_in_id_0 = r_766_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_15_io_in_id_1 = r_766_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_14_15_io_in_last_0 = r_1022_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_15_io_in_last_1 = r_1022_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_14_15_io_in_valid_0 = r_510_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_14_15_io_in_valid_1 = r_510_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_0_clock = clock;
  assign mesh_15_0_io_in_a_0 = r_240_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_0_io_in_a_1 = r_240_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_0_io_in_b_0 = pipe_b_15_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_b_1 = pipe_b_15_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_d_0 = pipe_b_271_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_d_1 = pipe_b_271_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_control_0_dataflow = mesh_15_0_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_control_0_propagate = mesh_15_0_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_control_0_shift = mesh_15_0_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_control_1_dataflow = mesh_15_0_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_control_1_propagate = mesh_15_0_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_control_1_shift = mesh_15_0_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_0_io_in_id_0 = r_527_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_0_io_in_id_1 = r_527_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_0_io_in_last_0 = r_783_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_0_io_in_last_1 = r_783_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_0_io_in_valid_0 = r_271_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_0_io_in_valid_1 = r_271_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_1_clock = clock;
  assign mesh_15_1_io_in_a_0 = r_241_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_1_io_in_a_1 = r_241_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_1_io_in_b_0 = pipe_b_31_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_b_1 = pipe_b_31_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_d_0 = pipe_b_287_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_d_1 = pipe_b_287_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_control_0_dataflow = mesh_15_1_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_control_0_propagate = mesh_15_1_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_control_0_shift = mesh_15_1_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_control_1_dataflow = mesh_15_1_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_control_1_propagate = mesh_15_1_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_control_1_shift = mesh_15_1_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_1_io_in_id_0 = r_543_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_1_io_in_id_1 = r_543_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_1_io_in_last_0 = r_799_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_1_io_in_last_1 = r_799_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_1_io_in_valid_0 = r_287_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_1_io_in_valid_1 = r_287_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_2_clock = clock;
  assign mesh_15_2_io_in_a_0 = r_242_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_2_io_in_a_1 = r_242_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_2_io_in_b_0 = pipe_b_47_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_b_1 = pipe_b_47_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_d_0 = pipe_b_303_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_d_1 = pipe_b_303_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_control_0_dataflow = mesh_15_2_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_control_0_propagate = mesh_15_2_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_control_0_shift = mesh_15_2_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_control_1_dataflow = mesh_15_2_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_control_1_propagate = mesh_15_2_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_control_1_shift = mesh_15_2_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_2_io_in_id_0 = r_559_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_2_io_in_id_1 = r_559_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_2_io_in_last_0 = r_815_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_2_io_in_last_1 = r_815_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_2_io_in_valid_0 = r_303_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_2_io_in_valid_1 = r_303_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_3_clock = clock;
  assign mesh_15_3_io_in_a_0 = r_243_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_3_io_in_a_1 = r_243_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_3_io_in_b_0 = pipe_b_63_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_b_1 = pipe_b_63_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_d_0 = pipe_b_319_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_d_1 = pipe_b_319_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_control_0_dataflow = mesh_15_3_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_control_0_propagate = mesh_15_3_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_control_0_shift = mesh_15_3_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_control_1_dataflow = mesh_15_3_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_control_1_propagate = mesh_15_3_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_control_1_shift = mesh_15_3_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_3_io_in_id_0 = r_575_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_3_io_in_id_1 = r_575_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_3_io_in_last_0 = r_831_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_3_io_in_last_1 = r_831_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_3_io_in_valid_0 = r_319_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_3_io_in_valid_1 = r_319_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_4_clock = clock;
  assign mesh_15_4_io_in_a_0 = r_244_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_4_io_in_a_1 = r_244_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_4_io_in_b_0 = pipe_b_79_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_b_1 = pipe_b_79_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_d_0 = pipe_b_335_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_d_1 = pipe_b_335_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_control_0_dataflow = mesh_15_4_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_control_0_propagate = mesh_15_4_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_control_0_shift = mesh_15_4_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_control_1_dataflow = mesh_15_4_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_control_1_propagate = mesh_15_4_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_control_1_shift = mesh_15_4_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_4_io_in_id_0 = r_591_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_4_io_in_id_1 = r_591_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_4_io_in_last_0 = r_847_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_4_io_in_last_1 = r_847_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_4_io_in_valid_0 = r_335_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_4_io_in_valid_1 = r_335_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_5_clock = clock;
  assign mesh_15_5_io_in_a_0 = r_245_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_5_io_in_a_1 = r_245_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_5_io_in_b_0 = pipe_b_95_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_b_1 = pipe_b_95_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_d_0 = pipe_b_351_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_d_1 = pipe_b_351_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_control_0_dataflow = mesh_15_5_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_control_0_propagate = mesh_15_5_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_control_0_shift = mesh_15_5_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_control_1_dataflow = mesh_15_5_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_control_1_propagate = mesh_15_5_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_control_1_shift = mesh_15_5_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_5_io_in_id_0 = r_607_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_5_io_in_id_1 = r_607_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_5_io_in_last_0 = r_863_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_5_io_in_last_1 = r_863_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_5_io_in_valid_0 = r_351_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_5_io_in_valid_1 = r_351_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_6_clock = clock;
  assign mesh_15_6_io_in_a_0 = r_246_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_6_io_in_a_1 = r_246_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_6_io_in_b_0 = pipe_b_111_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_b_1 = pipe_b_111_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_d_0 = pipe_b_367_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_d_1 = pipe_b_367_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_control_0_dataflow = mesh_15_6_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_control_0_propagate = mesh_15_6_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_control_0_shift = mesh_15_6_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_control_1_dataflow = mesh_15_6_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_control_1_propagate = mesh_15_6_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_control_1_shift = mesh_15_6_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_6_io_in_id_0 = r_623_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_6_io_in_id_1 = r_623_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_6_io_in_last_0 = r_879_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_6_io_in_last_1 = r_879_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_6_io_in_valid_0 = r_367_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_6_io_in_valid_1 = r_367_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_7_clock = clock;
  assign mesh_15_7_io_in_a_0 = r_247_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_7_io_in_a_1 = r_247_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_7_io_in_b_0 = pipe_b_127_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_b_1 = pipe_b_127_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_d_0 = pipe_b_383_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_d_1 = pipe_b_383_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_control_0_dataflow = mesh_15_7_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_control_0_propagate = mesh_15_7_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_control_0_shift = mesh_15_7_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_control_1_dataflow = mesh_15_7_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_control_1_propagate = mesh_15_7_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_control_1_shift = mesh_15_7_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_7_io_in_id_0 = r_639_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_7_io_in_id_1 = r_639_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_7_io_in_last_0 = r_895_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_7_io_in_last_1 = r_895_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_7_io_in_valid_0 = r_383_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_7_io_in_valid_1 = r_383_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_8_clock = clock;
  assign mesh_15_8_io_in_a_0 = r_248_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_8_io_in_a_1 = r_248_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_8_io_in_b_0 = pipe_b_143_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_b_1 = pipe_b_143_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_d_0 = pipe_b_399_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_d_1 = pipe_b_399_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_control_0_dataflow = mesh_15_8_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_control_0_propagate = mesh_15_8_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_control_0_shift = mesh_15_8_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_control_1_dataflow = mesh_15_8_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_control_1_propagate = mesh_15_8_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_control_1_shift = mesh_15_8_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_8_io_in_id_0 = r_655_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_8_io_in_id_1 = r_655_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_8_io_in_last_0 = r_911_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_8_io_in_last_1 = r_911_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_8_io_in_valid_0 = r_399_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_8_io_in_valid_1 = r_399_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_9_clock = clock;
  assign mesh_15_9_io_in_a_0 = r_249_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_9_io_in_a_1 = r_249_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_9_io_in_b_0 = pipe_b_159_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_b_1 = pipe_b_159_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_d_0 = pipe_b_415_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_d_1 = pipe_b_415_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_control_0_dataflow = mesh_15_9_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_control_0_propagate = mesh_15_9_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_control_0_shift = mesh_15_9_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_control_1_dataflow = mesh_15_9_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_control_1_propagate = mesh_15_9_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_control_1_shift = mesh_15_9_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_9_io_in_id_0 = r_671_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_9_io_in_id_1 = r_671_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_9_io_in_last_0 = r_927_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_9_io_in_last_1 = r_927_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_9_io_in_valid_0 = r_415_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_9_io_in_valid_1 = r_415_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_10_clock = clock;
  assign mesh_15_10_io_in_a_0 = r_250_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_10_io_in_a_1 = r_250_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_10_io_in_b_0 = pipe_b_175_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_b_1 = pipe_b_175_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_d_0 = pipe_b_431_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_d_1 = pipe_b_431_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_control_0_dataflow = mesh_15_10_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_control_0_propagate = mesh_15_10_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_control_0_shift = mesh_15_10_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_control_1_dataflow = mesh_15_10_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_control_1_propagate = mesh_15_10_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_control_1_shift = mesh_15_10_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_10_io_in_id_0 = r_687_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_10_io_in_id_1 = r_687_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_10_io_in_last_0 = r_943_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_10_io_in_last_1 = r_943_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_10_io_in_valid_0 = r_431_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_10_io_in_valid_1 = r_431_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_11_clock = clock;
  assign mesh_15_11_io_in_a_0 = r_251_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_11_io_in_a_1 = r_251_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_11_io_in_b_0 = pipe_b_191_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_b_1 = pipe_b_191_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_d_0 = pipe_b_447_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_d_1 = pipe_b_447_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_control_0_dataflow = mesh_15_11_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_control_0_propagate = mesh_15_11_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_control_0_shift = mesh_15_11_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_control_1_dataflow = mesh_15_11_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_control_1_propagate = mesh_15_11_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_control_1_shift = mesh_15_11_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_11_io_in_id_0 = r_703_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_11_io_in_id_1 = r_703_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_11_io_in_last_0 = r_959_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_11_io_in_last_1 = r_959_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_11_io_in_valid_0 = r_447_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_11_io_in_valid_1 = r_447_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_12_clock = clock;
  assign mesh_15_12_io_in_a_0 = r_252_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_12_io_in_a_1 = r_252_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_12_io_in_b_0 = pipe_b_207_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_b_1 = pipe_b_207_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_d_0 = pipe_b_463_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_d_1 = pipe_b_463_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_control_0_dataflow = mesh_15_12_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_control_0_propagate = mesh_15_12_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_control_0_shift = mesh_15_12_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_control_1_dataflow = mesh_15_12_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_control_1_propagate = mesh_15_12_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_control_1_shift = mesh_15_12_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_12_io_in_id_0 = r_719_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_12_io_in_id_1 = r_719_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_12_io_in_last_0 = r_975_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_12_io_in_last_1 = r_975_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_12_io_in_valid_0 = r_463_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_12_io_in_valid_1 = r_463_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_13_clock = clock;
  assign mesh_15_13_io_in_a_0 = r_253_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_13_io_in_a_1 = r_253_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_13_io_in_b_0 = pipe_b_223_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_b_1 = pipe_b_223_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_d_0 = pipe_b_479_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_d_1 = pipe_b_479_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_control_0_dataflow = mesh_15_13_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_control_0_propagate = mesh_15_13_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_control_0_shift = mesh_15_13_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_control_1_dataflow = mesh_15_13_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_control_1_propagate = mesh_15_13_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_control_1_shift = mesh_15_13_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_13_io_in_id_0 = r_735_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_13_io_in_id_1 = r_735_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_13_io_in_last_0 = r_991_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_13_io_in_last_1 = r_991_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_13_io_in_valid_0 = r_479_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_13_io_in_valid_1 = r_479_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_14_clock = clock;
  assign mesh_15_14_io_in_a_0 = r_254_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_14_io_in_a_1 = r_254_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_14_io_in_b_0 = pipe_b_239_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_b_1 = pipe_b_239_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_d_0 = pipe_b_495_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_d_1 = pipe_b_495_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_control_0_dataflow = mesh_15_14_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_control_0_propagate = mesh_15_14_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_control_0_shift = mesh_15_14_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_control_1_dataflow = mesh_15_14_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_control_1_propagate = mesh_15_14_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_control_1_shift = mesh_15_14_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_14_io_in_id_0 = r_751_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_14_io_in_id_1 = r_751_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_14_io_in_last_0 = r_1007_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_14_io_in_last_1 = r_1007_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_14_io_in_valid_0 = r_495_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_14_io_in_valid_1 = r_495_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_15_clock = clock;
  assign mesh_15_15_io_in_a_0 = r_255_0; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_15_io_in_a_1 = r_255_1; // @[src/main/scala/gemmini/Mesh.scala 53:22]
  assign mesh_15_15_io_in_b_0 = pipe_b_255_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_b_1 = pipe_b_255_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_d_0 = pipe_b_511_0; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_d_1 = pipe_b_511_1; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_control_0_dataflow = mesh_15_15_io_in_control_0_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_control_0_propagate = mesh_15_15_io_in_control_0_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_control_0_shift = mesh_15_15_io_in_control_0_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_control_1_dataflow = mesh_15_15_io_in_control_1_dataflow_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_control_1_propagate = mesh_15_15_io_in_control_1_propagate_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_control_1_shift = mesh_15_15_io_in_control_1_shift_pipe_b; // @[src/main/scala/chisel3/util/Valid.scala 128:21 130:16]
  assign mesh_15_15_io_in_id_0 = r_767_0; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_15_io_in_id_1 = r_767_1; // @[src/main/scala/gemmini/Mesh.scala 103:23]
  assign mesh_15_15_io_in_last_0 = r_1023_0; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_15_io_in_last_1 = r_1023_1; // @[src/main/scala/gemmini/Mesh.scala 112:25]
  assign mesh_15_15_io_in_valid_0 = r_511_0; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  assign mesh_15_15_io_in_valid_1 = r_511_1; // @[src/main/scala/gemmini/Mesh.scala 94:26]
  always @(posedge clock) begin
    r__0 <= io_in_a_0_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r__1 <= io_in_a_0_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_1_0 <= mesh_0_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_1_1 <= mesh_0_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_2_0 <= mesh_0_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_2_1 <= mesh_0_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_3_0 <= mesh_0_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_3_1 <= mesh_0_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_4_0 <= mesh_0_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_4_1 <= mesh_0_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_5_0 <= mesh_0_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_5_1 <= mesh_0_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_6_0 <= mesh_0_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_6_1 <= mesh_0_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_7_0 <= mesh_0_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_7_1 <= mesh_0_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_8_0 <= mesh_0_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_8_1 <= mesh_0_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_9_0 <= mesh_0_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_9_1 <= mesh_0_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_10_0 <= mesh_0_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_10_1 <= mesh_0_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_11_0 <= mesh_0_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_11_1 <= mesh_0_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_12_0 <= mesh_0_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_12_1 <= mesh_0_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_13_0 <= mesh_0_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_13_1 <= mesh_0_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_14_0 <= mesh_0_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_14_1 <= mesh_0_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_15_0 <= mesh_0_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_15_1 <= mesh_0_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_16_0 <= io_in_a_1_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_16_1 <= io_in_a_1_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_17_0 <= mesh_1_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_17_1 <= mesh_1_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_18_0 <= mesh_1_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_18_1 <= mesh_1_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_19_0 <= mesh_1_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_19_1 <= mesh_1_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_20_0 <= mesh_1_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_20_1 <= mesh_1_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_21_0 <= mesh_1_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_21_1 <= mesh_1_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_22_0 <= mesh_1_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_22_1 <= mesh_1_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_23_0 <= mesh_1_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_23_1 <= mesh_1_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_24_0 <= mesh_1_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_24_1 <= mesh_1_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_25_0 <= mesh_1_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_25_1 <= mesh_1_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_26_0 <= mesh_1_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_26_1 <= mesh_1_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_27_0 <= mesh_1_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_27_1 <= mesh_1_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_28_0 <= mesh_1_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_28_1 <= mesh_1_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_29_0 <= mesh_1_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_29_1 <= mesh_1_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_30_0 <= mesh_1_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_30_1 <= mesh_1_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_31_0 <= mesh_1_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_31_1 <= mesh_1_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_32_0 <= io_in_a_2_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_32_1 <= io_in_a_2_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_33_0 <= mesh_2_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_33_1 <= mesh_2_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_34_0 <= mesh_2_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_34_1 <= mesh_2_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_35_0 <= mesh_2_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_35_1 <= mesh_2_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_36_0 <= mesh_2_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_36_1 <= mesh_2_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_37_0 <= mesh_2_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_37_1 <= mesh_2_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_38_0 <= mesh_2_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_38_1 <= mesh_2_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_39_0 <= mesh_2_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_39_1 <= mesh_2_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_40_0 <= mesh_2_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_40_1 <= mesh_2_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_41_0 <= mesh_2_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_41_1 <= mesh_2_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_42_0 <= mesh_2_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_42_1 <= mesh_2_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_43_0 <= mesh_2_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_43_1 <= mesh_2_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_44_0 <= mesh_2_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_44_1 <= mesh_2_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_45_0 <= mesh_2_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_45_1 <= mesh_2_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_46_0 <= mesh_2_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_46_1 <= mesh_2_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_47_0 <= mesh_2_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_47_1 <= mesh_2_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_48_0 <= io_in_a_3_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_48_1 <= io_in_a_3_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_49_0 <= mesh_3_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_49_1 <= mesh_3_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_50_0 <= mesh_3_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_50_1 <= mesh_3_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_51_0 <= mesh_3_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_51_1 <= mesh_3_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_52_0 <= mesh_3_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_52_1 <= mesh_3_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_53_0 <= mesh_3_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_53_1 <= mesh_3_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_54_0 <= mesh_3_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_54_1 <= mesh_3_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_55_0 <= mesh_3_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_55_1 <= mesh_3_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_56_0 <= mesh_3_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_56_1 <= mesh_3_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_57_0 <= mesh_3_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_57_1 <= mesh_3_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_58_0 <= mesh_3_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_58_1 <= mesh_3_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_59_0 <= mesh_3_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_59_1 <= mesh_3_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_60_0 <= mesh_3_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_60_1 <= mesh_3_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_61_0 <= mesh_3_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_61_1 <= mesh_3_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_62_0 <= mesh_3_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_62_1 <= mesh_3_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_63_0 <= mesh_3_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_63_1 <= mesh_3_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_64_0 <= io_in_a_4_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_64_1 <= io_in_a_4_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_65_0 <= mesh_4_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_65_1 <= mesh_4_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_66_0 <= mesh_4_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_66_1 <= mesh_4_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_67_0 <= mesh_4_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_67_1 <= mesh_4_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_68_0 <= mesh_4_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_68_1 <= mesh_4_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_69_0 <= mesh_4_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_69_1 <= mesh_4_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_70_0 <= mesh_4_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_70_1 <= mesh_4_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_71_0 <= mesh_4_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_71_1 <= mesh_4_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_72_0 <= mesh_4_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_72_1 <= mesh_4_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_73_0 <= mesh_4_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_73_1 <= mesh_4_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_74_0 <= mesh_4_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_74_1 <= mesh_4_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_75_0 <= mesh_4_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_75_1 <= mesh_4_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_76_0 <= mesh_4_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_76_1 <= mesh_4_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_77_0 <= mesh_4_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_77_1 <= mesh_4_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_78_0 <= mesh_4_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_78_1 <= mesh_4_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_79_0 <= mesh_4_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_79_1 <= mesh_4_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_80_0 <= io_in_a_5_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_80_1 <= io_in_a_5_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_81_0 <= mesh_5_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_81_1 <= mesh_5_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_82_0 <= mesh_5_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_82_1 <= mesh_5_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_83_0 <= mesh_5_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_83_1 <= mesh_5_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_84_0 <= mesh_5_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_84_1 <= mesh_5_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_85_0 <= mesh_5_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_85_1 <= mesh_5_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_86_0 <= mesh_5_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_86_1 <= mesh_5_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_87_0 <= mesh_5_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_87_1 <= mesh_5_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_88_0 <= mesh_5_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_88_1 <= mesh_5_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_89_0 <= mesh_5_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_89_1 <= mesh_5_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_90_0 <= mesh_5_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_90_1 <= mesh_5_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_91_0 <= mesh_5_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_91_1 <= mesh_5_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_92_0 <= mesh_5_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_92_1 <= mesh_5_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_93_0 <= mesh_5_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_93_1 <= mesh_5_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_94_0 <= mesh_5_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_94_1 <= mesh_5_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_95_0 <= mesh_5_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_95_1 <= mesh_5_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_96_0 <= io_in_a_6_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_96_1 <= io_in_a_6_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_97_0 <= mesh_6_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_97_1 <= mesh_6_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_98_0 <= mesh_6_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_98_1 <= mesh_6_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_99_0 <= mesh_6_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_99_1 <= mesh_6_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_100_0 <= mesh_6_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_100_1 <= mesh_6_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_101_0 <= mesh_6_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_101_1 <= mesh_6_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_102_0 <= mesh_6_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_102_1 <= mesh_6_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_103_0 <= mesh_6_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_103_1 <= mesh_6_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_104_0 <= mesh_6_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_104_1 <= mesh_6_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_105_0 <= mesh_6_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_105_1 <= mesh_6_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_106_0 <= mesh_6_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_106_1 <= mesh_6_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_107_0 <= mesh_6_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_107_1 <= mesh_6_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_108_0 <= mesh_6_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_108_1 <= mesh_6_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_109_0 <= mesh_6_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_109_1 <= mesh_6_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_110_0 <= mesh_6_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_110_1 <= mesh_6_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_111_0 <= mesh_6_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_111_1 <= mesh_6_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_112_0 <= io_in_a_7_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_112_1 <= io_in_a_7_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_113_0 <= mesh_7_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_113_1 <= mesh_7_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_114_0 <= mesh_7_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_114_1 <= mesh_7_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_115_0 <= mesh_7_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_115_1 <= mesh_7_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_116_0 <= mesh_7_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_116_1 <= mesh_7_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_117_0 <= mesh_7_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_117_1 <= mesh_7_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_118_0 <= mesh_7_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_118_1 <= mesh_7_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_119_0 <= mesh_7_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_119_1 <= mesh_7_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_120_0 <= mesh_7_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_120_1 <= mesh_7_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_121_0 <= mesh_7_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_121_1 <= mesh_7_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_122_0 <= mesh_7_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_122_1 <= mesh_7_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_123_0 <= mesh_7_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_123_1 <= mesh_7_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_124_0 <= mesh_7_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_124_1 <= mesh_7_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_125_0 <= mesh_7_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_125_1 <= mesh_7_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_126_0 <= mesh_7_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_126_1 <= mesh_7_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_127_0 <= mesh_7_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_127_1 <= mesh_7_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_128_0 <= io_in_a_8_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_128_1 <= io_in_a_8_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_129_0 <= mesh_8_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_129_1 <= mesh_8_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_130_0 <= mesh_8_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_130_1 <= mesh_8_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_131_0 <= mesh_8_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_131_1 <= mesh_8_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_132_0 <= mesh_8_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_132_1 <= mesh_8_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_133_0 <= mesh_8_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_133_1 <= mesh_8_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_134_0 <= mesh_8_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_134_1 <= mesh_8_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_135_0 <= mesh_8_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_135_1 <= mesh_8_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_136_0 <= mesh_8_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_136_1 <= mesh_8_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_137_0 <= mesh_8_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_137_1 <= mesh_8_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_138_0 <= mesh_8_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_138_1 <= mesh_8_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_139_0 <= mesh_8_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_139_1 <= mesh_8_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_140_0 <= mesh_8_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_140_1 <= mesh_8_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_141_0 <= mesh_8_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_141_1 <= mesh_8_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_142_0 <= mesh_8_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_142_1 <= mesh_8_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_143_0 <= mesh_8_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_143_1 <= mesh_8_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_144_0 <= io_in_a_9_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_144_1 <= io_in_a_9_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_145_0 <= mesh_9_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_145_1 <= mesh_9_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_146_0 <= mesh_9_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_146_1 <= mesh_9_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_147_0 <= mesh_9_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_147_1 <= mesh_9_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_148_0 <= mesh_9_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_148_1 <= mesh_9_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_149_0 <= mesh_9_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_149_1 <= mesh_9_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_150_0 <= mesh_9_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_150_1 <= mesh_9_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_151_0 <= mesh_9_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_151_1 <= mesh_9_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_152_0 <= mesh_9_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_152_1 <= mesh_9_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_153_0 <= mesh_9_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_153_1 <= mesh_9_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_154_0 <= mesh_9_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_154_1 <= mesh_9_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_155_0 <= mesh_9_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_155_1 <= mesh_9_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_156_0 <= mesh_9_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_156_1 <= mesh_9_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_157_0 <= mesh_9_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_157_1 <= mesh_9_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_158_0 <= mesh_9_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_158_1 <= mesh_9_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_159_0 <= mesh_9_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_159_1 <= mesh_9_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_160_0 <= io_in_a_10_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_160_1 <= io_in_a_10_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_161_0 <= mesh_10_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_161_1 <= mesh_10_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_162_0 <= mesh_10_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_162_1 <= mesh_10_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_163_0 <= mesh_10_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_163_1 <= mesh_10_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_164_0 <= mesh_10_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_164_1 <= mesh_10_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_165_0 <= mesh_10_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_165_1 <= mesh_10_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_166_0 <= mesh_10_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_166_1 <= mesh_10_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_167_0 <= mesh_10_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_167_1 <= mesh_10_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_168_0 <= mesh_10_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_168_1 <= mesh_10_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_169_0 <= mesh_10_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_169_1 <= mesh_10_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_170_0 <= mesh_10_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_170_1 <= mesh_10_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_171_0 <= mesh_10_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_171_1 <= mesh_10_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_172_0 <= mesh_10_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_172_1 <= mesh_10_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_173_0 <= mesh_10_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_173_1 <= mesh_10_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_174_0 <= mesh_10_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_174_1 <= mesh_10_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_175_0 <= mesh_10_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_175_1 <= mesh_10_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_176_0 <= io_in_a_11_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_176_1 <= io_in_a_11_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_177_0 <= mesh_11_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_177_1 <= mesh_11_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_178_0 <= mesh_11_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_178_1 <= mesh_11_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_179_0 <= mesh_11_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_179_1 <= mesh_11_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_180_0 <= mesh_11_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_180_1 <= mesh_11_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_181_0 <= mesh_11_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_181_1 <= mesh_11_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_182_0 <= mesh_11_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_182_1 <= mesh_11_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_183_0 <= mesh_11_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_183_1 <= mesh_11_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_184_0 <= mesh_11_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_184_1 <= mesh_11_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_185_0 <= mesh_11_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_185_1 <= mesh_11_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_186_0 <= mesh_11_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_186_1 <= mesh_11_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_187_0 <= mesh_11_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_187_1 <= mesh_11_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_188_0 <= mesh_11_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_188_1 <= mesh_11_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_189_0 <= mesh_11_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_189_1 <= mesh_11_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_190_0 <= mesh_11_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_190_1 <= mesh_11_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_191_0 <= mesh_11_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_191_1 <= mesh_11_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_192_0 <= io_in_a_12_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_192_1 <= io_in_a_12_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_193_0 <= mesh_12_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_193_1 <= mesh_12_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_194_0 <= mesh_12_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_194_1 <= mesh_12_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_195_0 <= mesh_12_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_195_1 <= mesh_12_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_196_0 <= mesh_12_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_196_1 <= mesh_12_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_197_0 <= mesh_12_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_197_1 <= mesh_12_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_198_0 <= mesh_12_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_198_1 <= mesh_12_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_199_0 <= mesh_12_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_199_1 <= mesh_12_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_200_0 <= mesh_12_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_200_1 <= mesh_12_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_201_0 <= mesh_12_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_201_1 <= mesh_12_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_202_0 <= mesh_12_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_202_1 <= mesh_12_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_203_0 <= mesh_12_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_203_1 <= mesh_12_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_204_0 <= mesh_12_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_204_1 <= mesh_12_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_205_0 <= mesh_12_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_205_1 <= mesh_12_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_206_0 <= mesh_12_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_206_1 <= mesh_12_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_207_0 <= mesh_12_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_207_1 <= mesh_12_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_208_0 <= io_in_a_13_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_208_1 <= io_in_a_13_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_209_0 <= mesh_13_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_209_1 <= mesh_13_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_210_0 <= mesh_13_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_210_1 <= mesh_13_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_211_0 <= mesh_13_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_211_1 <= mesh_13_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_212_0 <= mesh_13_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_212_1 <= mesh_13_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_213_0 <= mesh_13_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_213_1 <= mesh_13_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_214_0 <= mesh_13_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_214_1 <= mesh_13_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_215_0 <= mesh_13_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_215_1 <= mesh_13_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_216_0 <= mesh_13_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_216_1 <= mesh_13_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_217_0 <= mesh_13_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_217_1 <= mesh_13_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_218_0 <= mesh_13_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_218_1 <= mesh_13_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_219_0 <= mesh_13_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_219_1 <= mesh_13_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_220_0 <= mesh_13_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_220_1 <= mesh_13_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_221_0 <= mesh_13_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_221_1 <= mesh_13_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_222_0 <= mesh_13_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_222_1 <= mesh_13_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_223_0 <= mesh_13_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_223_1 <= mesh_13_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_224_0 <= io_in_a_14_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_224_1 <= io_in_a_14_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_225_0 <= mesh_14_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_225_1 <= mesh_14_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_226_0 <= mesh_14_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_226_1 <= mesh_14_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_227_0 <= mesh_14_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_227_1 <= mesh_14_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_228_0 <= mesh_14_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_228_1 <= mesh_14_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_229_0 <= mesh_14_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_229_1 <= mesh_14_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_230_0 <= mesh_14_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_230_1 <= mesh_14_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_231_0 <= mesh_14_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_231_1 <= mesh_14_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_232_0 <= mesh_14_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_232_1 <= mesh_14_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_233_0 <= mesh_14_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_233_1 <= mesh_14_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_234_0 <= mesh_14_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_234_1 <= mesh_14_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_235_0 <= mesh_14_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_235_1 <= mesh_14_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_236_0 <= mesh_14_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_236_1 <= mesh_14_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_237_0 <= mesh_14_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_237_1 <= mesh_14_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_238_0 <= mesh_14_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_238_1 <= mesh_14_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_239_0 <= mesh_14_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_239_1 <= mesh_14_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_240_0 <= io_in_a_15_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_240_1 <= io_in_a_15_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_241_0 <= mesh_15_0_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_241_1 <= mesh_15_0_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_242_0 <= mesh_15_1_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_242_1 <= mesh_15_1_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_243_0 <= mesh_15_2_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_243_1 <= mesh_15_2_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_244_0 <= mesh_15_3_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_244_1 <= mesh_15_3_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_245_0 <= mesh_15_4_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_245_1 <= mesh_15_4_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_246_0 <= mesh_15_5_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_246_1 <= mesh_15_5_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_247_0 <= mesh_15_6_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_247_1 <= mesh_15_6_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_248_0 <= mesh_15_7_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_248_1 <= mesh_15_7_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_249_0 <= mesh_15_8_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_249_1 <= mesh_15_8_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_250_0 <= mesh_15_9_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_250_1 <= mesh_15_9_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_251_0 <= mesh_15_10_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_251_1 <= mesh_15_10_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_252_0 <= mesh_15_11_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_252_1 <= mesh_15_11_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_253_0 <= mesh_15_12_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_253_1 <= mesh_15_12_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_254_0 <= mesh_15_13_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_254_1 <= mesh_15_13_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_255_0 <= mesh_15_14_io_out_a_0; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    r_255_1 <= mesh_15_14_io_out_a_1; // @[src/main/scala/gemmini/Mesh.scala 53:{38,38,38}]
    if (io_in_valid_0_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b__0 <= io_in_b_0_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b__1 <= io_in_b_0_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_1_0 <= mesh_0_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_1_1 <= mesh_0_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_2_0 <= mesh_1_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_2_1 <= mesh_1_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_3_0 <= mesh_2_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_3_1 <= mesh_2_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_4_0 <= mesh_3_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_4_1 <= mesh_3_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_5_0 <= mesh_4_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_5_1 <= mesh_4_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_6_0 <= mesh_5_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_6_1 <= mesh_5_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_7_0 <= mesh_6_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_7_1 <= mesh_6_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_8_0 <= mesh_7_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_8_1 <= mesh_7_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_9_0 <= mesh_8_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_9_1 <= mesh_8_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_10_0 <= mesh_9_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_10_1 <= mesh_9_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_11_0 <= mesh_10_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_11_1 <= mesh_10_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_12_0 <= mesh_11_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_12_1 <= mesh_11_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_13_0 <= mesh_12_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_13_1 <= mesh_12_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_14_0 <= mesh_13_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_14_1 <= mesh_13_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_15_0 <= mesh_14_0_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_15_1 <= mesh_14_0_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_16_0 <= io_in_b_1_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_16_1 <= io_in_b_1_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_17_0 <= mesh_0_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_17_1 <= mesh_0_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_18_0 <= mesh_1_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_18_1 <= mesh_1_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_19_0 <= mesh_2_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_19_1 <= mesh_2_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_20_0 <= mesh_3_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_20_1 <= mesh_3_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_21_0 <= mesh_4_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_21_1 <= mesh_4_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_22_0 <= mesh_5_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_22_1 <= mesh_5_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_23_0 <= mesh_6_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_23_1 <= mesh_6_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_24_0 <= mesh_7_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_24_1 <= mesh_7_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_25_0 <= mesh_8_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_25_1 <= mesh_8_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_26_0 <= mesh_9_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_26_1 <= mesh_9_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_27_0 <= mesh_10_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_27_1 <= mesh_10_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_28_0 <= mesh_11_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_28_1 <= mesh_11_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_29_0 <= mesh_12_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_29_1 <= mesh_12_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_30_0 <= mesh_13_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_30_1 <= mesh_13_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_31_0 <= mesh_14_1_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_31_1 <= mesh_14_1_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_32_0 <= io_in_b_2_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_32_1 <= io_in_b_2_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_33_0 <= mesh_0_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_33_1 <= mesh_0_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_34_0 <= mesh_1_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_34_1 <= mesh_1_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_35_0 <= mesh_2_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_35_1 <= mesh_2_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_36_0 <= mesh_3_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_36_1 <= mesh_3_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_37_0 <= mesh_4_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_37_1 <= mesh_4_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_38_0 <= mesh_5_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_38_1 <= mesh_5_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_39_0 <= mesh_6_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_39_1 <= mesh_6_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_40_0 <= mesh_7_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_40_1 <= mesh_7_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_41_0 <= mesh_8_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_41_1 <= mesh_8_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_42_0 <= mesh_9_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_42_1 <= mesh_9_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_43_0 <= mesh_10_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_43_1 <= mesh_10_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_44_0 <= mesh_11_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_44_1 <= mesh_11_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_45_0 <= mesh_12_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_45_1 <= mesh_12_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_46_0 <= mesh_13_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_46_1 <= mesh_13_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_47_0 <= mesh_14_2_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_47_1 <= mesh_14_2_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_48_0 <= io_in_b_3_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_48_1 <= io_in_b_3_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_49_0 <= mesh_0_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_49_1 <= mesh_0_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_50_0 <= mesh_1_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_50_1 <= mesh_1_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_51_0 <= mesh_2_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_51_1 <= mesh_2_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_52_0 <= mesh_3_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_52_1 <= mesh_3_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_53_0 <= mesh_4_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_53_1 <= mesh_4_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_54_0 <= mesh_5_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_54_1 <= mesh_5_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_55_0 <= mesh_6_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_55_1 <= mesh_6_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_56_0 <= mesh_7_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_56_1 <= mesh_7_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_57_0 <= mesh_8_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_57_1 <= mesh_8_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_58_0 <= mesh_9_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_58_1 <= mesh_9_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_59_0 <= mesh_10_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_59_1 <= mesh_10_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_60_0 <= mesh_11_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_60_1 <= mesh_11_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_61_0 <= mesh_12_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_61_1 <= mesh_12_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_62_0 <= mesh_13_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_62_1 <= mesh_13_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_63_0 <= mesh_14_3_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_63_1 <= mesh_14_3_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_64_0 <= io_in_b_4_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_64_1 <= io_in_b_4_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_65_0 <= mesh_0_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_65_1 <= mesh_0_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_66_0 <= mesh_1_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_66_1 <= mesh_1_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_67_0 <= mesh_2_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_67_1 <= mesh_2_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_68_0 <= mesh_3_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_68_1 <= mesh_3_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_69_0 <= mesh_4_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_69_1 <= mesh_4_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_70_0 <= mesh_5_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_70_1 <= mesh_5_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_71_0 <= mesh_6_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_71_1 <= mesh_6_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_72_0 <= mesh_7_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_72_1 <= mesh_7_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_73_0 <= mesh_8_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_73_1 <= mesh_8_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_74_0 <= mesh_9_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_74_1 <= mesh_9_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_75_0 <= mesh_10_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_75_1 <= mesh_10_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_76_0 <= mesh_11_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_76_1 <= mesh_11_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_77_0 <= mesh_12_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_77_1 <= mesh_12_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_78_0 <= mesh_13_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_78_1 <= mesh_13_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_79_0 <= mesh_14_4_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_79_1 <= mesh_14_4_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_80_0 <= io_in_b_5_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_80_1 <= io_in_b_5_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_81_0 <= mesh_0_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_81_1 <= mesh_0_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_82_0 <= mesh_1_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_82_1 <= mesh_1_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_83_0 <= mesh_2_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_83_1 <= mesh_2_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_84_0 <= mesh_3_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_84_1 <= mesh_3_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_85_0 <= mesh_4_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_85_1 <= mesh_4_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_86_0 <= mesh_5_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_86_1 <= mesh_5_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_87_0 <= mesh_6_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_87_1 <= mesh_6_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_88_0 <= mesh_7_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_88_1 <= mesh_7_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_89_0 <= mesh_8_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_89_1 <= mesh_8_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_90_0 <= mesh_9_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_90_1 <= mesh_9_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_91_0 <= mesh_10_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_91_1 <= mesh_10_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_92_0 <= mesh_11_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_92_1 <= mesh_11_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_93_0 <= mesh_12_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_93_1 <= mesh_12_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_94_0 <= mesh_13_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_94_1 <= mesh_13_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_95_0 <= mesh_14_5_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_95_1 <= mesh_14_5_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_96_0 <= io_in_b_6_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_96_1 <= io_in_b_6_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_97_0 <= mesh_0_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_97_1 <= mesh_0_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_98_0 <= mesh_1_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_98_1 <= mesh_1_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_99_0 <= mesh_2_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_99_1 <= mesh_2_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_100_0 <= mesh_3_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_100_1 <= mesh_3_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_101_0 <= mesh_4_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_101_1 <= mesh_4_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_102_0 <= mesh_5_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_102_1 <= mesh_5_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_103_0 <= mesh_6_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_103_1 <= mesh_6_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_104_0 <= mesh_7_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_104_1 <= mesh_7_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_105_0 <= mesh_8_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_105_1 <= mesh_8_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_106_0 <= mesh_9_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_106_1 <= mesh_9_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_107_0 <= mesh_10_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_107_1 <= mesh_10_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_108_0 <= mesh_11_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_108_1 <= mesh_11_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_109_0 <= mesh_12_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_109_1 <= mesh_12_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_110_0 <= mesh_13_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_110_1 <= mesh_13_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_111_0 <= mesh_14_6_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_111_1 <= mesh_14_6_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_112_0 <= io_in_b_7_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_112_1 <= io_in_b_7_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_113_0 <= mesh_0_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_113_1 <= mesh_0_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_114_0 <= mesh_1_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_114_1 <= mesh_1_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_115_0 <= mesh_2_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_115_1 <= mesh_2_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_116_0 <= mesh_3_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_116_1 <= mesh_3_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_117_0 <= mesh_4_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_117_1 <= mesh_4_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_118_0 <= mesh_5_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_118_1 <= mesh_5_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_119_0 <= mesh_6_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_119_1 <= mesh_6_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_120_0 <= mesh_7_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_120_1 <= mesh_7_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_121_0 <= mesh_8_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_121_1 <= mesh_8_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_122_0 <= mesh_9_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_122_1 <= mesh_9_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_123_0 <= mesh_10_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_123_1 <= mesh_10_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_124_0 <= mesh_11_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_124_1 <= mesh_11_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_125_0 <= mesh_12_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_125_1 <= mesh_12_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_126_0 <= mesh_13_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_126_1 <= mesh_13_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_127_0 <= mesh_14_7_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_127_1 <= mesh_14_7_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_128_0 <= io_in_b_8_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_128_1 <= io_in_b_8_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_129_0 <= mesh_0_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_129_1 <= mesh_0_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_130_0 <= mesh_1_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_130_1 <= mesh_1_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_131_0 <= mesh_2_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_131_1 <= mesh_2_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_132_0 <= mesh_3_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_132_1 <= mesh_3_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_133_0 <= mesh_4_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_133_1 <= mesh_4_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_134_0 <= mesh_5_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_134_1 <= mesh_5_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_135_0 <= mesh_6_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_135_1 <= mesh_6_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_136_0 <= mesh_7_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_136_1 <= mesh_7_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_137_0 <= mesh_8_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_137_1 <= mesh_8_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_138_0 <= mesh_9_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_138_1 <= mesh_9_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_139_0 <= mesh_10_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_139_1 <= mesh_10_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_140_0 <= mesh_11_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_140_1 <= mesh_11_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_141_0 <= mesh_12_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_141_1 <= mesh_12_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_142_0 <= mesh_13_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_142_1 <= mesh_13_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_143_0 <= mesh_14_8_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_143_1 <= mesh_14_8_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_144_0 <= io_in_b_9_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_144_1 <= io_in_b_9_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_145_0 <= mesh_0_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_145_1 <= mesh_0_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_146_0 <= mesh_1_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_146_1 <= mesh_1_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_147_0 <= mesh_2_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_147_1 <= mesh_2_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_148_0 <= mesh_3_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_148_1 <= mesh_3_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_149_0 <= mesh_4_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_149_1 <= mesh_4_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_150_0 <= mesh_5_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_150_1 <= mesh_5_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_151_0 <= mesh_6_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_151_1 <= mesh_6_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_152_0 <= mesh_7_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_152_1 <= mesh_7_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_153_0 <= mesh_8_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_153_1 <= mesh_8_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_154_0 <= mesh_9_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_154_1 <= mesh_9_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_155_0 <= mesh_10_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_155_1 <= mesh_10_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_156_0 <= mesh_11_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_156_1 <= mesh_11_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_157_0 <= mesh_12_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_157_1 <= mesh_12_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_158_0 <= mesh_13_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_158_1 <= mesh_13_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_159_0 <= mesh_14_9_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_159_1 <= mesh_14_9_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_160_0 <= io_in_b_10_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_160_1 <= io_in_b_10_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_161_0 <= mesh_0_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_161_1 <= mesh_0_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_162_0 <= mesh_1_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_162_1 <= mesh_1_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_163_0 <= mesh_2_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_163_1 <= mesh_2_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_164_0 <= mesh_3_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_164_1 <= mesh_3_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_165_0 <= mesh_4_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_165_1 <= mesh_4_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_166_0 <= mesh_5_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_166_1 <= mesh_5_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_167_0 <= mesh_6_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_167_1 <= mesh_6_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_168_0 <= mesh_7_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_168_1 <= mesh_7_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_169_0 <= mesh_8_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_169_1 <= mesh_8_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_170_0 <= mesh_9_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_170_1 <= mesh_9_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_171_0 <= mesh_10_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_171_1 <= mesh_10_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_172_0 <= mesh_11_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_172_1 <= mesh_11_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_173_0 <= mesh_12_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_173_1 <= mesh_12_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_174_0 <= mesh_13_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_174_1 <= mesh_13_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_175_0 <= mesh_14_10_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_175_1 <= mesh_14_10_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_176_0 <= io_in_b_11_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_176_1 <= io_in_b_11_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_177_0 <= mesh_0_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_177_1 <= mesh_0_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_178_0 <= mesh_1_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_178_1 <= mesh_1_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_179_0 <= mesh_2_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_179_1 <= mesh_2_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_180_0 <= mesh_3_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_180_1 <= mesh_3_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_181_0 <= mesh_4_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_181_1 <= mesh_4_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_182_0 <= mesh_5_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_182_1 <= mesh_5_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_183_0 <= mesh_6_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_183_1 <= mesh_6_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_184_0 <= mesh_7_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_184_1 <= mesh_7_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_185_0 <= mesh_8_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_185_1 <= mesh_8_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_186_0 <= mesh_9_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_186_1 <= mesh_9_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_187_0 <= mesh_10_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_187_1 <= mesh_10_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_188_0 <= mesh_11_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_188_1 <= mesh_11_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_189_0 <= mesh_12_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_189_1 <= mesh_12_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_190_0 <= mesh_13_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_190_1 <= mesh_13_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_191_0 <= mesh_14_11_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_191_1 <= mesh_14_11_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_192_0 <= io_in_b_12_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_192_1 <= io_in_b_12_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_193_0 <= mesh_0_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_193_1 <= mesh_0_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_194_0 <= mesh_1_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_194_1 <= mesh_1_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_195_0 <= mesh_2_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_195_1 <= mesh_2_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_196_0 <= mesh_3_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_196_1 <= mesh_3_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_197_0 <= mesh_4_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_197_1 <= mesh_4_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_198_0 <= mesh_5_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_198_1 <= mesh_5_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_199_0 <= mesh_6_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_199_1 <= mesh_6_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_200_0 <= mesh_7_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_200_1 <= mesh_7_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_201_0 <= mesh_8_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_201_1 <= mesh_8_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_202_0 <= mesh_9_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_202_1 <= mesh_9_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_203_0 <= mesh_10_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_203_1 <= mesh_10_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_204_0 <= mesh_11_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_204_1 <= mesh_11_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_205_0 <= mesh_12_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_205_1 <= mesh_12_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_206_0 <= mesh_13_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_206_1 <= mesh_13_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_207_0 <= mesh_14_12_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_207_1 <= mesh_14_12_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_208_0 <= io_in_b_13_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_208_1 <= io_in_b_13_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_209_0 <= mesh_0_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_209_1 <= mesh_0_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_210_0 <= mesh_1_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_210_1 <= mesh_1_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_211_0 <= mesh_2_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_211_1 <= mesh_2_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_212_0 <= mesh_3_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_212_1 <= mesh_3_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_213_0 <= mesh_4_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_213_1 <= mesh_4_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_214_0 <= mesh_5_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_214_1 <= mesh_5_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_215_0 <= mesh_6_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_215_1 <= mesh_6_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_216_0 <= mesh_7_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_216_1 <= mesh_7_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_217_0 <= mesh_8_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_217_1 <= mesh_8_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_218_0 <= mesh_9_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_218_1 <= mesh_9_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_219_0 <= mesh_10_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_219_1 <= mesh_10_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_220_0 <= mesh_11_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_220_1 <= mesh_11_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_221_0 <= mesh_12_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_221_1 <= mesh_12_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_222_0 <= mesh_13_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_222_1 <= mesh_13_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_223_0 <= mesh_14_13_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_223_1 <= mesh_14_13_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_224_0 <= io_in_b_14_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_224_1 <= io_in_b_14_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_225_0 <= mesh_0_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_225_1 <= mesh_0_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_226_0 <= mesh_1_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_226_1 <= mesh_1_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_227_0 <= mesh_2_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_227_1 <= mesh_2_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_228_0 <= mesh_3_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_228_1 <= mesh_3_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_229_0 <= mesh_4_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_229_1 <= mesh_4_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_230_0 <= mesh_5_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_230_1 <= mesh_5_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_231_0 <= mesh_6_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_231_1 <= mesh_6_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_232_0 <= mesh_7_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_232_1 <= mesh_7_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_233_0 <= mesh_8_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_233_1 <= mesh_8_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_234_0 <= mesh_9_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_234_1 <= mesh_9_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_235_0 <= mesh_10_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_235_1 <= mesh_10_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_236_0 <= mesh_11_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_236_1 <= mesh_11_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_237_0 <= mesh_12_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_237_1 <= mesh_12_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_238_0 <= mesh_13_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_238_1 <= mesh_13_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_239_0 <= mesh_14_14_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_239_1 <= mesh_14_14_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_240_0 <= io_in_b_15_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_240_1 <= io_in_b_15_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_241_0 <= mesh_0_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_241_1 <= mesh_0_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_242_0 <= mesh_1_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_242_1 <= mesh_1_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_243_0 <= mesh_2_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_243_1 <= mesh_2_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_244_0 <= mesh_3_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_244_1 <= mesh_3_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_245_0 <= mesh_4_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_245_1 <= mesh_4_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_246_0 <= mesh_5_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_246_1 <= mesh_5_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_247_0 <= mesh_6_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_247_1 <= mesh_6_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_248_0 <= mesh_7_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_248_1 <= mesh_7_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_249_0 <= mesh_8_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_249_1 <= mesh_8_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_250_0 <= mesh_9_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_250_1 <= mesh_9_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_251_0 <= mesh_10_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_251_1 <= mesh_10_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_252_0 <= mesh_11_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_252_1 <= mesh_11_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_253_0 <= mesh_12_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_253_1 <= mesh_12_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_254_0 <= mesh_13_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_254_1 <= mesh_13_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_255_0 <= mesh_14_15_io_out_b_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_255_1 <= mesh_14_15_io_out_b_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_256_0 <= io_in_d_0_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_256_1 <= io_in_d_0_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_257_0 <= mesh_0_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_257_1 <= mesh_0_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_258_0 <= mesh_1_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_258_1 <= mesh_1_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_259_0 <= mesh_2_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_259_1 <= mesh_2_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_260_0 <= mesh_3_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_260_1 <= mesh_3_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_261_0 <= mesh_4_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_261_1 <= mesh_4_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_262_0 <= mesh_5_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_262_1 <= mesh_5_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_263_0 <= mesh_6_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_263_1 <= mesh_6_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_264_0 <= mesh_7_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_264_1 <= mesh_7_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_265_0 <= mesh_8_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_265_1 <= mesh_8_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_266_0 <= mesh_9_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_266_1 <= mesh_9_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_267_0 <= mesh_10_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_267_1 <= mesh_10_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_268_0 <= mesh_11_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_268_1 <= mesh_11_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_269_0 <= mesh_12_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_269_1 <= mesh_12_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_270_0 <= mesh_13_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_270_1 <= mesh_13_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_271_0 <= mesh_14_0_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_271_1 <= mesh_14_0_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_272_0 <= io_in_d_1_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_272_1 <= io_in_d_1_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_273_0 <= mesh_0_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_273_1 <= mesh_0_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_274_0 <= mesh_1_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_274_1 <= mesh_1_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_275_0 <= mesh_2_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_275_1 <= mesh_2_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_276_0 <= mesh_3_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_276_1 <= mesh_3_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_277_0 <= mesh_4_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_277_1 <= mesh_4_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_278_0 <= mesh_5_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_278_1 <= mesh_5_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_279_0 <= mesh_6_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_279_1 <= mesh_6_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_280_0 <= mesh_7_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_280_1 <= mesh_7_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_281_0 <= mesh_8_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_281_1 <= mesh_8_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_282_0 <= mesh_9_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_282_1 <= mesh_9_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_283_0 <= mesh_10_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_283_1 <= mesh_10_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_284_0 <= mesh_11_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_284_1 <= mesh_11_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_285_0 <= mesh_12_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_285_1 <= mesh_12_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_286_0 <= mesh_13_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_286_1 <= mesh_13_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_287_0 <= mesh_14_1_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_287_1 <= mesh_14_1_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_288_0 <= io_in_d_2_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_288_1 <= io_in_d_2_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_289_0 <= mesh_0_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_289_1 <= mesh_0_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_290_0 <= mesh_1_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_290_1 <= mesh_1_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_291_0 <= mesh_2_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_291_1 <= mesh_2_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_292_0 <= mesh_3_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_292_1 <= mesh_3_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_293_0 <= mesh_4_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_293_1 <= mesh_4_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_294_0 <= mesh_5_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_294_1 <= mesh_5_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_295_0 <= mesh_6_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_295_1 <= mesh_6_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_296_0 <= mesh_7_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_296_1 <= mesh_7_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_297_0 <= mesh_8_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_297_1 <= mesh_8_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_298_0 <= mesh_9_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_298_1 <= mesh_9_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_299_0 <= mesh_10_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_299_1 <= mesh_10_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_300_0 <= mesh_11_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_300_1 <= mesh_11_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_301_0 <= mesh_12_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_301_1 <= mesh_12_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_302_0 <= mesh_13_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_302_1 <= mesh_13_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_303_0 <= mesh_14_2_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_303_1 <= mesh_14_2_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_304_0 <= io_in_d_3_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_304_1 <= io_in_d_3_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_305_0 <= mesh_0_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_305_1 <= mesh_0_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_306_0 <= mesh_1_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_306_1 <= mesh_1_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_307_0 <= mesh_2_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_307_1 <= mesh_2_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_308_0 <= mesh_3_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_308_1 <= mesh_3_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_309_0 <= mesh_4_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_309_1 <= mesh_4_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_310_0 <= mesh_5_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_310_1 <= mesh_5_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_311_0 <= mesh_6_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_311_1 <= mesh_6_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_312_0 <= mesh_7_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_312_1 <= mesh_7_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_313_0 <= mesh_8_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_313_1 <= mesh_8_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_314_0 <= mesh_9_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_314_1 <= mesh_9_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_315_0 <= mesh_10_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_315_1 <= mesh_10_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_316_0 <= mesh_11_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_316_1 <= mesh_11_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_317_0 <= mesh_12_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_317_1 <= mesh_12_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_318_0 <= mesh_13_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_318_1 <= mesh_13_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_319_0 <= mesh_14_3_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_319_1 <= mesh_14_3_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_320_0 <= io_in_d_4_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_320_1 <= io_in_d_4_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_321_0 <= mesh_0_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_321_1 <= mesh_0_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_322_0 <= mesh_1_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_322_1 <= mesh_1_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_323_0 <= mesh_2_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_323_1 <= mesh_2_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_324_0 <= mesh_3_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_324_1 <= mesh_3_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_325_0 <= mesh_4_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_325_1 <= mesh_4_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_326_0 <= mesh_5_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_326_1 <= mesh_5_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_327_0 <= mesh_6_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_327_1 <= mesh_6_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_328_0 <= mesh_7_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_328_1 <= mesh_7_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_329_0 <= mesh_8_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_329_1 <= mesh_8_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_330_0 <= mesh_9_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_330_1 <= mesh_9_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_331_0 <= mesh_10_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_331_1 <= mesh_10_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_332_0 <= mesh_11_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_332_1 <= mesh_11_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_333_0 <= mesh_12_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_333_1 <= mesh_12_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_334_0 <= mesh_13_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_334_1 <= mesh_13_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_335_0 <= mesh_14_4_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_335_1 <= mesh_14_4_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_336_0 <= io_in_d_5_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_336_1 <= io_in_d_5_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_337_0 <= mesh_0_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_337_1 <= mesh_0_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_338_0 <= mesh_1_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_338_1 <= mesh_1_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_339_0 <= mesh_2_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_339_1 <= mesh_2_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_340_0 <= mesh_3_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_340_1 <= mesh_3_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_341_0 <= mesh_4_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_341_1 <= mesh_4_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_342_0 <= mesh_5_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_342_1 <= mesh_5_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_343_0 <= mesh_6_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_343_1 <= mesh_6_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_344_0 <= mesh_7_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_344_1 <= mesh_7_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_345_0 <= mesh_8_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_345_1 <= mesh_8_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_346_0 <= mesh_9_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_346_1 <= mesh_9_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_347_0 <= mesh_10_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_347_1 <= mesh_10_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_348_0 <= mesh_11_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_348_1 <= mesh_11_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_349_0 <= mesh_12_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_349_1 <= mesh_12_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_350_0 <= mesh_13_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_350_1 <= mesh_13_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_351_0 <= mesh_14_5_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_351_1 <= mesh_14_5_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_352_0 <= io_in_d_6_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_352_1 <= io_in_d_6_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_353_0 <= mesh_0_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_353_1 <= mesh_0_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_354_0 <= mesh_1_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_354_1 <= mesh_1_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_355_0 <= mesh_2_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_355_1 <= mesh_2_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_356_0 <= mesh_3_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_356_1 <= mesh_3_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_357_0 <= mesh_4_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_357_1 <= mesh_4_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_358_0 <= mesh_5_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_358_1 <= mesh_5_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_359_0 <= mesh_6_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_359_1 <= mesh_6_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_360_0 <= mesh_7_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_360_1 <= mesh_7_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_361_0 <= mesh_8_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_361_1 <= mesh_8_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_362_0 <= mesh_9_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_362_1 <= mesh_9_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_363_0 <= mesh_10_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_363_1 <= mesh_10_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_364_0 <= mesh_11_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_364_1 <= mesh_11_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_365_0 <= mesh_12_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_365_1 <= mesh_12_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_366_0 <= mesh_13_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_366_1 <= mesh_13_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_367_0 <= mesh_14_6_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_367_1 <= mesh_14_6_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_368_0 <= io_in_d_7_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_368_1 <= io_in_d_7_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_369_0 <= mesh_0_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_369_1 <= mesh_0_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_370_0 <= mesh_1_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_370_1 <= mesh_1_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_371_0 <= mesh_2_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_371_1 <= mesh_2_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_372_0 <= mesh_3_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_372_1 <= mesh_3_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_373_0 <= mesh_4_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_373_1 <= mesh_4_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_374_0 <= mesh_5_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_374_1 <= mesh_5_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_375_0 <= mesh_6_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_375_1 <= mesh_6_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_376_0 <= mesh_7_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_376_1 <= mesh_7_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_377_0 <= mesh_8_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_377_1 <= mesh_8_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_378_0 <= mesh_9_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_378_1 <= mesh_9_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_379_0 <= mesh_10_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_379_1 <= mesh_10_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_380_0 <= mesh_11_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_380_1 <= mesh_11_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_381_0 <= mesh_12_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_381_1 <= mesh_12_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_382_0 <= mesh_13_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_382_1 <= mesh_13_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_383_0 <= mesh_14_7_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_383_1 <= mesh_14_7_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_384_0 <= io_in_d_8_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_384_1 <= io_in_d_8_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_385_0 <= mesh_0_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_385_1 <= mesh_0_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_386_0 <= mesh_1_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_386_1 <= mesh_1_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_387_0 <= mesh_2_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_387_1 <= mesh_2_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_388_0 <= mesh_3_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_388_1 <= mesh_3_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_389_0 <= mesh_4_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_389_1 <= mesh_4_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_390_0 <= mesh_5_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_390_1 <= mesh_5_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_391_0 <= mesh_6_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_391_1 <= mesh_6_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_392_0 <= mesh_7_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_392_1 <= mesh_7_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_393_0 <= mesh_8_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_393_1 <= mesh_8_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_394_0 <= mesh_9_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_394_1 <= mesh_9_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_395_0 <= mesh_10_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_395_1 <= mesh_10_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_396_0 <= mesh_11_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_396_1 <= mesh_11_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_397_0 <= mesh_12_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_397_1 <= mesh_12_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_398_0 <= mesh_13_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_398_1 <= mesh_13_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_399_0 <= mesh_14_8_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_399_1 <= mesh_14_8_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_400_0 <= io_in_d_9_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_400_1 <= io_in_d_9_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_401_0 <= mesh_0_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_401_1 <= mesh_0_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_402_0 <= mesh_1_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_402_1 <= mesh_1_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_403_0 <= mesh_2_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_403_1 <= mesh_2_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_404_0 <= mesh_3_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_404_1 <= mesh_3_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_405_0 <= mesh_4_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_405_1 <= mesh_4_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_406_0 <= mesh_5_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_406_1 <= mesh_5_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_407_0 <= mesh_6_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_407_1 <= mesh_6_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_408_0 <= mesh_7_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_408_1 <= mesh_7_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_409_0 <= mesh_8_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_409_1 <= mesh_8_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_410_0 <= mesh_9_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_410_1 <= mesh_9_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_411_0 <= mesh_10_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_411_1 <= mesh_10_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_412_0 <= mesh_11_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_412_1 <= mesh_11_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_413_0 <= mesh_12_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_413_1 <= mesh_12_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_414_0 <= mesh_13_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_414_1 <= mesh_13_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_415_0 <= mesh_14_9_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_415_1 <= mesh_14_9_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_416_0 <= io_in_d_10_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_416_1 <= io_in_d_10_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_417_0 <= mesh_0_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_417_1 <= mesh_0_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_418_0 <= mesh_1_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_418_1 <= mesh_1_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_419_0 <= mesh_2_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_419_1 <= mesh_2_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_420_0 <= mesh_3_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_420_1 <= mesh_3_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_421_0 <= mesh_4_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_421_1 <= mesh_4_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_422_0 <= mesh_5_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_422_1 <= mesh_5_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_423_0 <= mesh_6_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_423_1 <= mesh_6_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_424_0 <= mesh_7_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_424_1 <= mesh_7_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_425_0 <= mesh_8_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_425_1 <= mesh_8_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_426_0 <= mesh_9_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_426_1 <= mesh_9_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_427_0 <= mesh_10_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_427_1 <= mesh_10_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_428_0 <= mesh_11_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_428_1 <= mesh_11_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_429_0 <= mesh_12_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_429_1 <= mesh_12_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_430_0 <= mesh_13_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_430_1 <= mesh_13_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_431_0 <= mesh_14_10_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_431_1 <= mesh_14_10_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_432_0 <= io_in_d_11_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_432_1 <= io_in_d_11_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_433_0 <= mesh_0_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_433_1 <= mesh_0_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_434_0 <= mesh_1_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_434_1 <= mesh_1_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_435_0 <= mesh_2_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_435_1 <= mesh_2_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_436_0 <= mesh_3_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_436_1 <= mesh_3_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_437_0 <= mesh_4_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_437_1 <= mesh_4_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_438_0 <= mesh_5_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_438_1 <= mesh_5_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_439_0 <= mesh_6_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_439_1 <= mesh_6_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_440_0 <= mesh_7_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_440_1 <= mesh_7_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_441_0 <= mesh_8_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_441_1 <= mesh_8_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_442_0 <= mesh_9_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_442_1 <= mesh_9_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_443_0 <= mesh_10_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_443_1 <= mesh_10_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_444_0 <= mesh_11_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_444_1 <= mesh_11_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_445_0 <= mesh_12_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_445_1 <= mesh_12_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_446_0 <= mesh_13_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_446_1 <= mesh_13_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_447_0 <= mesh_14_11_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_447_1 <= mesh_14_11_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_448_0 <= io_in_d_12_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_448_1 <= io_in_d_12_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_449_0 <= mesh_0_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_449_1 <= mesh_0_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_450_0 <= mesh_1_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_450_1 <= mesh_1_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_451_0 <= mesh_2_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_451_1 <= mesh_2_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_452_0 <= mesh_3_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_452_1 <= mesh_3_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_453_0 <= mesh_4_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_453_1 <= mesh_4_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_454_0 <= mesh_5_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_454_1 <= mesh_5_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_455_0 <= mesh_6_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_455_1 <= mesh_6_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_456_0 <= mesh_7_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_456_1 <= mesh_7_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_457_0 <= mesh_8_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_457_1 <= mesh_8_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_458_0 <= mesh_9_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_458_1 <= mesh_9_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_459_0 <= mesh_10_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_459_1 <= mesh_10_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_460_0 <= mesh_11_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_460_1 <= mesh_11_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_461_0 <= mesh_12_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_461_1 <= mesh_12_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_462_0 <= mesh_13_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_462_1 <= mesh_13_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_463_0 <= mesh_14_12_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_463_1 <= mesh_14_12_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_464_0 <= io_in_d_13_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_464_1 <= io_in_d_13_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_465_0 <= mesh_0_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_465_1 <= mesh_0_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_466_0 <= mesh_1_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_466_1 <= mesh_1_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_467_0 <= mesh_2_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_467_1 <= mesh_2_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_468_0 <= mesh_3_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_468_1 <= mesh_3_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_469_0 <= mesh_4_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_469_1 <= mesh_4_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_470_0 <= mesh_5_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_470_1 <= mesh_5_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_471_0 <= mesh_6_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_471_1 <= mesh_6_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_472_0 <= mesh_7_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_472_1 <= mesh_7_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_473_0 <= mesh_8_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_473_1 <= mesh_8_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_474_0 <= mesh_9_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_474_1 <= mesh_9_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_475_0 <= mesh_10_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_475_1 <= mesh_10_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_476_0 <= mesh_11_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_476_1 <= mesh_11_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_477_0 <= mesh_12_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_477_1 <= mesh_12_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_478_0 <= mesh_13_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_478_1 <= mesh_13_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_479_0 <= mesh_14_13_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_479_1 <= mesh_14_13_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_480_0 <= io_in_d_14_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_480_1 <= io_in_d_14_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_481_0 <= mesh_0_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_481_1 <= mesh_0_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_482_0 <= mesh_1_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_482_1 <= mesh_1_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_483_0 <= mesh_2_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_483_1 <= mesh_2_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_484_0 <= mesh_3_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_484_1 <= mesh_3_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_485_0 <= mesh_4_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_485_1 <= mesh_4_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_486_0 <= mesh_5_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_486_1 <= mesh_5_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_487_0 <= mesh_6_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_487_1 <= mesh_6_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_488_0 <= mesh_7_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_488_1 <= mesh_7_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_489_0 <= mesh_8_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_489_1 <= mesh_8_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_490_0 <= mesh_9_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_490_1 <= mesh_9_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_491_0 <= mesh_10_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_491_1 <= mesh_10_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_492_0 <= mesh_11_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_492_1 <= mesh_11_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_493_0 <= mesh_12_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_493_1 <= mesh_12_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_494_0 <= mesh_13_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_494_1 <= mesh_13_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_495_0 <= mesh_14_14_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_495_1 <= mesh_14_14_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_496_0 <= io_in_d_15_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_496_1 <= io_in_d_15_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_497_0 <= mesh_0_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_497_1 <= mesh_0_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_498_0 <= mesh_1_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_498_1 <= mesh_1_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_499_0 <= mesh_2_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_499_1 <= mesh_2_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_500_0 <= mesh_3_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_500_1 <= mesh_3_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_501_0 <= mesh_4_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_501_1 <= mesh_4_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_502_0 <= mesh_5_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_502_1 <= mesh_5_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_503_0 <= mesh_6_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_503_1 <= mesh_6_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_504_0 <= mesh_7_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_504_1 <= mesh_7_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_505_0 <= mesh_8_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_505_1 <= mesh_8_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_506_0 <= mesh_9_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_506_1 <= mesh_9_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_507_0 <= mesh_10_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_507_1 <= mesh_10_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_508_0 <= mesh_11_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_508_1 <= mesh_11_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_509_0 <= mesh_12_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_509_1 <= mesh_12_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_510_0 <= mesh_13_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_510_1 <= mesh_13_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_511_0 <= mesh_14_15_io_out_c_0; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      pipe_b_511_1 <= mesh_14_15_io_out_c_1; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_0_io_in_control_0_shift_pipe_b <= io_in_control_0_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_0_io_in_control_0_dataflow_pipe_b <= io_in_control_0_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_0_io_in_control_0_propagate_pipe_b <= io_in_control_0_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_0_io_in_control_1_shift_pipe_b <= io_in_control_0_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_0_io_in_control_1_dataflow_pipe_b <= io_in_control_0_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_0_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_0_io_in_control_1_propagate_pipe_b <= io_in_control_0_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_0_io_in_control_0_shift_pipe_b <= mesh_0_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_0_io_in_control_0_dataflow_pipe_b <= mesh_0_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_0_io_in_control_0_propagate_pipe_b <= mesh_0_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_0_io_in_control_1_shift_pipe_b <= mesh_0_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_0_io_in_control_1_dataflow_pipe_b <= mesh_0_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_0_io_in_control_1_propagate_pipe_b <= mesh_0_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_0_io_in_control_0_shift_pipe_b <= mesh_1_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_0_io_in_control_0_dataflow_pipe_b <= mesh_1_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_0_io_in_control_0_propagate_pipe_b <= mesh_1_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_0_io_in_control_1_shift_pipe_b <= mesh_1_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_0_io_in_control_1_dataflow_pipe_b <= mesh_1_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_0_io_in_control_1_propagate_pipe_b <= mesh_1_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_0_io_in_control_0_shift_pipe_b <= mesh_2_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_0_io_in_control_0_dataflow_pipe_b <= mesh_2_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_0_io_in_control_0_propagate_pipe_b <= mesh_2_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_0_io_in_control_1_shift_pipe_b <= mesh_2_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_0_io_in_control_1_dataflow_pipe_b <= mesh_2_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_0_io_in_control_1_propagate_pipe_b <= mesh_2_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_0_io_in_control_0_shift_pipe_b <= mesh_3_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_0_io_in_control_0_dataflow_pipe_b <= mesh_3_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_0_io_in_control_0_propagate_pipe_b <= mesh_3_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_0_io_in_control_1_shift_pipe_b <= mesh_3_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_0_io_in_control_1_dataflow_pipe_b <= mesh_3_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_0_io_in_control_1_propagate_pipe_b <= mesh_3_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_0_io_in_control_0_shift_pipe_b <= mesh_4_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_0_io_in_control_0_dataflow_pipe_b <= mesh_4_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_0_io_in_control_0_propagate_pipe_b <= mesh_4_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_0_io_in_control_1_shift_pipe_b <= mesh_4_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_0_io_in_control_1_dataflow_pipe_b <= mesh_4_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_0_io_in_control_1_propagate_pipe_b <= mesh_4_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_0_io_in_control_0_shift_pipe_b <= mesh_5_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_0_io_in_control_0_dataflow_pipe_b <= mesh_5_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_0_io_in_control_0_propagate_pipe_b <= mesh_5_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_0_io_in_control_1_shift_pipe_b <= mesh_5_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_0_io_in_control_1_dataflow_pipe_b <= mesh_5_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_0_io_in_control_1_propagate_pipe_b <= mesh_5_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_0_io_in_control_0_shift_pipe_b <= mesh_6_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_0_io_in_control_0_dataflow_pipe_b <= mesh_6_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_0_io_in_control_0_propagate_pipe_b <= mesh_6_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_0_io_in_control_1_shift_pipe_b <= mesh_6_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_0_io_in_control_1_dataflow_pipe_b <= mesh_6_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_0_io_in_control_1_propagate_pipe_b <= mesh_6_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_0_io_in_control_0_shift_pipe_b <= mesh_7_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_0_io_in_control_0_dataflow_pipe_b <= mesh_7_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_0_io_in_control_0_propagate_pipe_b <= mesh_7_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_0_io_in_control_1_shift_pipe_b <= mesh_7_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_0_io_in_control_1_dataflow_pipe_b <= mesh_7_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_0_io_in_control_1_propagate_pipe_b <= mesh_7_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_0_io_in_control_0_shift_pipe_b <= mesh_8_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_0_io_in_control_0_dataflow_pipe_b <= mesh_8_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_0_io_in_control_0_propagate_pipe_b <= mesh_8_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_0_io_in_control_1_shift_pipe_b <= mesh_8_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_0_io_in_control_1_dataflow_pipe_b <= mesh_8_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_0_io_in_control_1_propagate_pipe_b <= mesh_8_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_0_io_in_control_0_shift_pipe_b <= mesh_9_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_0_io_in_control_0_dataflow_pipe_b <= mesh_9_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_0_io_in_control_0_propagate_pipe_b <= mesh_9_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_0_io_in_control_1_shift_pipe_b <= mesh_9_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_0_io_in_control_1_dataflow_pipe_b <= mesh_9_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_0_io_in_control_1_propagate_pipe_b <= mesh_9_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_0_io_in_control_0_shift_pipe_b <= mesh_10_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_0_io_in_control_0_dataflow_pipe_b <= mesh_10_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_0_io_in_control_0_propagate_pipe_b <= mesh_10_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_0_io_in_control_1_shift_pipe_b <= mesh_10_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_0_io_in_control_1_dataflow_pipe_b <= mesh_10_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_0_io_in_control_1_propagate_pipe_b <= mesh_10_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_0_io_in_control_0_shift_pipe_b <= mesh_11_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_0_io_in_control_0_dataflow_pipe_b <= mesh_11_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_0_io_in_control_0_propagate_pipe_b <= mesh_11_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_0_io_in_control_1_shift_pipe_b <= mesh_11_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_0_io_in_control_1_dataflow_pipe_b <= mesh_11_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_0_io_in_control_1_propagate_pipe_b <= mesh_11_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_0_io_in_control_0_shift_pipe_b <= mesh_12_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_0_io_in_control_0_dataflow_pipe_b <= mesh_12_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_0_io_in_control_0_propagate_pipe_b <= mesh_12_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_0_io_in_control_1_shift_pipe_b <= mesh_12_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_0_io_in_control_1_dataflow_pipe_b <= mesh_12_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_0_io_in_control_1_propagate_pipe_b <= mesh_12_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_0_io_in_control_0_shift_pipe_b <= mesh_13_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_0_io_in_control_0_dataflow_pipe_b <= mesh_13_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_0_io_in_control_0_propagate_pipe_b <= mesh_13_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_0_io_in_control_1_shift_pipe_b <= mesh_13_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_0_io_in_control_1_dataflow_pipe_b <= mesh_13_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_0_io_in_control_1_propagate_pipe_b <= mesh_13_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_0_io_in_control_0_shift_pipe_b <= mesh_14_0_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_0_io_in_control_0_dataflow_pipe_b <= mesh_14_0_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_0_io_in_control_0_propagate_pipe_b <= mesh_14_0_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_0_io_in_control_1_shift_pipe_b <= mesh_14_0_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_0_io_in_control_1_dataflow_pipe_b <= mesh_14_0_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_0_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_0_io_in_control_1_propagate_pipe_b <= mesh_14_0_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_1_io_in_control_0_shift_pipe_b <= io_in_control_1_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_1_io_in_control_0_dataflow_pipe_b <= io_in_control_1_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_1_io_in_control_0_propagate_pipe_b <= io_in_control_1_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_1_io_in_control_1_shift_pipe_b <= io_in_control_1_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_1_io_in_control_1_dataflow_pipe_b <= io_in_control_1_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_1_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_1_io_in_control_1_propagate_pipe_b <= io_in_control_1_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_1_io_in_control_0_shift_pipe_b <= mesh_0_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_1_io_in_control_0_dataflow_pipe_b <= mesh_0_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_1_io_in_control_0_propagate_pipe_b <= mesh_0_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_1_io_in_control_1_shift_pipe_b <= mesh_0_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_1_io_in_control_1_dataflow_pipe_b <= mesh_0_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_1_io_in_control_1_propagate_pipe_b <= mesh_0_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_1_io_in_control_0_shift_pipe_b <= mesh_1_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_1_io_in_control_0_dataflow_pipe_b <= mesh_1_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_1_io_in_control_0_propagate_pipe_b <= mesh_1_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_1_io_in_control_1_shift_pipe_b <= mesh_1_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_1_io_in_control_1_dataflow_pipe_b <= mesh_1_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_1_io_in_control_1_propagate_pipe_b <= mesh_1_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_1_io_in_control_0_shift_pipe_b <= mesh_2_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_1_io_in_control_0_dataflow_pipe_b <= mesh_2_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_1_io_in_control_0_propagate_pipe_b <= mesh_2_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_1_io_in_control_1_shift_pipe_b <= mesh_2_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_1_io_in_control_1_dataflow_pipe_b <= mesh_2_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_1_io_in_control_1_propagate_pipe_b <= mesh_2_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_1_io_in_control_0_shift_pipe_b <= mesh_3_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_1_io_in_control_0_dataflow_pipe_b <= mesh_3_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_1_io_in_control_0_propagate_pipe_b <= mesh_3_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_1_io_in_control_1_shift_pipe_b <= mesh_3_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_1_io_in_control_1_dataflow_pipe_b <= mesh_3_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_1_io_in_control_1_propagate_pipe_b <= mesh_3_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_1_io_in_control_0_shift_pipe_b <= mesh_4_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_1_io_in_control_0_dataflow_pipe_b <= mesh_4_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_1_io_in_control_0_propagate_pipe_b <= mesh_4_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_1_io_in_control_1_shift_pipe_b <= mesh_4_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_1_io_in_control_1_dataflow_pipe_b <= mesh_4_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_1_io_in_control_1_propagate_pipe_b <= mesh_4_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_1_io_in_control_0_shift_pipe_b <= mesh_5_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_1_io_in_control_0_dataflow_pipe_b <= mesh_5_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_1_io_in_control_0_propagate_pipe_b <= mesh_5_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_1_io_in_control_1_shift_pipe_b <= mesh_5_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_1_io_in_control_1_dataflow_pipe_b <= mesh_5_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_1_io_in_control_1_propagate_pipe_b <= mesh_5_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_1_io_in_control_0_shift_pipe_b <= mesh_6_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_1_io_in_control_0_dataflow_pipe_b <= mesh_6_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_1_io_in_control_0_propagate_pipe_b <= mesh_6_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_1_io_in_control_1_shift_pipe_b <= mesh_6_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_1_io_in_control_1_dataflow_pipe_b <= mesh_6_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_1_io_in_control_1_propagate_pipe_b <= mesh_6_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_1_io_in_control_0_shift_pipe_b <= mesh_7_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_1_io_in_control_0_dataflow_pipe_b <= mesh_7_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_1_io_in_control_0_propagate_pipe_b <= mesh_7_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_1_io_in_control_1_shift_pipe_b <= mesh_7_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_1_io_in_control_1_dataflow_pipe_b <= mesh_7_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_1_io_in_control_1_propagate_pipe_b <= mesh_7_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_1_io_in_control_0_shift_pipe_b <= mesh_8_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_1_io_in_control_0_dataflow_pipe_b <= mesh_8_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_1_io_in_control_0_propagate_pipe_b <= mesh_8_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_1_io_in_control_1_shift_pipe_b <= mesh_8_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_1_io_in_control_1_dataflow_pipe_b <= mesh_8_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_1_io_in_control_1_propagate_pipe_b <= mesh_8_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_1_io_in_control_0_shift_pipe_b <= mesh_9_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_1_io_in_control_0_dataflow_pipe_b <= mesh_9_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_1_io_in_control_0_propagate_pipe_b <= mesh_9_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_1_io_in_control_1_shift_pipe_b <= mesh_9_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_1_io_in_control_1_dataflow_pipe_b <= mesh_9_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_1_io_in_control_1_propagate_pipe_b <= mesh_9_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_1_io_in_control_0_shift_pipe_b <= mesh_10_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_1_io_in_control_0_dataflow_pipe_b <= mesh_10_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_1_io_in_control_0_propagate_pipe_b <= mesh_10_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_1_io_in_control_1_shift_pipe_b <= mesh_10_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_1_io_in_control_1_dataflow_pipe_b <= mesh_10_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_1_io_in_control_1_propagate_pipe_b <= mesh_10_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_1_io_in_control_0_shift_pipe_b <= mesh_11_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_1_io_in_control_0_dataflow_pipe_b <= mesh_11_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_1_io_in_control_0_propagate_pipe_b <= mesh_11_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_1_io_in_control_1_shift_pipe_b <= mesh_11_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_1_io_in_control_1_dataflow_pipe_b <= mesh_11_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_1_io_in_control_1_propagate_pipe_b <= mesh_11_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_1_io_in_control_0_shift_pipe_b <= mesh_12_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_1_io_in_control_0_dataflow_pipe_b <= mesh_12_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_1_io_in_control_0_propagate_pipe_b <= mesh_12_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_1_io_in_control_1_shift_pipe_b <= mesh_12_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_1_io_in_control_1_dataflow_pipe_b <= mesh_12_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_1_io_in_control_1_propagate_pipe_b <= mesh_12_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_1_io_in_control_0_shift_pipe_b <= mesh_13_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_1_io_in_control_0_dataflow_pipe_b <= mesh_13_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_1_io_in_control_0_propagate_pipe_b <= mesh_13_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_1_io_in_control_1_shift_pipe_b <= mesh_13_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_1_io_in_control_1_dataflow_pipe_b <= mesh_13_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_1_io_in_control_1_propagate_pipe_b <= mesh_13_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_1_io_in_control_0_shift_pipe_b <= mesh_14_1_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_1_io_in_control_0_dataflow_pipe_b <= mesh_14_1_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_1_io_in_control_0_propagate_pipe_b <= mesh_14_1_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_1_io_in_control_1_shift_pipe_b <= mesh_14_1_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_1_io_in_control_1_dataflow_pipe_b <= mesh_14_1_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_1_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_1_io_in_control_1_propagate_pipe_b <= mesh_14_1_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_2_io_in_control_0_shift_pipe_b <= io_in_control_2_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_2_io_in_control_0_dataflow_pipe_b <= io_in_control_2_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_2_io_in_control_0_propagate_pipe_b <= io_in_control_2_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_2_io_in_control_1_shift_pipe_b <= io_in_control_2_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_2_io_in_control_1_dataflow_pipe_b <= io_in_control_2_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_2_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_2_io_in_control_1_propagate_pipe_b <= io_in_control_2_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_2_io_in_control_0_shift_pipe_b <= mesh_0_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_2_io_in_control_0_dataflow_pipe_b <= mesh_0_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_2_io_in_control_0_propagate_pipe_b <= mesh_0_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_2_io_in_control_1_shift_pipe_b <= mesh_0_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_2_io_in_control_1_dataflow_pipe_b <= mesh_0_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_2_io_in_control_1_propagate_pipe_b <= mesh_0_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_2_io_in_control_0_shift_pipe_b <= mesh_1_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_2_io_in_control_0_dataflow_pipe_b <= mesh_1_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_2_io_in_control_0_propagate_pipe_b <= mesh_1_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_2_io_in_control_1_shift_pipe_b <= mesh_1_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_2_io_in_control_1_dataflow_pipe_b <= mesh_1_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_2_io_in_control_1_propagate_pipe_b <= mesh_1_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_2_io_in_control_0_shift_pipe_b <= mesh_2_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_2_io_in_control_0_dataflow_pipe_b <= mesh_2_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_2_io_in_control_0_propagate_pipe_b <= mesh_2_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_2_io_in_control_1_shift_pipe_b <= mesh_2_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_2_io_in_control_1_dataflow_pipe_b <= mesh_2_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_2_io_in_control_1_propagate_pipe_b <= mesh_2_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_2_io_in_control_0_shift_pipe_b <= mesh_3_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_2_io_in_control_0_dataflow_pipe_b <= mesh_3_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_2_io_in_control_0_propagate_pipe_b <= mesh_3_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_2_io_in_control_1_shift_pipe_b <= mesh_3_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_2_io_in_control_1_dataflow_pipe_b <= mesh_3_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_2_io_in_control_1_propagate_pipe_b <= mesh_3_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_2_io_in_control_0_shift_pipe_b <= mesh_4_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_2_io_in_control_0_dataflow_pipe_b <= mesh_4_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_2_io_in_control_0_propagate_pipe_b <= mesh_4_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_2_io_in_control_1_shift_pipe_b <= mesh_4_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_2_io_in_control_1_dataflow_pipe_b <= mesh_4_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_2_io_in_control_1_propagate_pipe_b <= mesh_4_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_2_io_in_control_0_shift_pipe_b <= mesh_5_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_2_io_in_control_0_dataflow_pipe_b <= mesh_5_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_2_io_in_control_0_propagate_pipe_b <= mesh_5_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_2_io_in_control_1_shift_pipe_b <= mesh_5_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_2_io_in_control_1_dataflow_pipe_b <= mesh_5_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_2_io_in_control_1_propagate_pipe_b <= mesh_5_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_2_io_in_control_0_shift_pipe_b <= mesh_6_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_2_io_in_control_0_dataflow_pipe_b <= mesh_6_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_2_io_in_control_0_propagate_pipe_b <= mesh_6_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_2_io_in_control_1_shift_pipe_b <= mesh_6_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_2_io_in_control_1_dataflow_pipe_b <= mesh_6_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_2_io_in_control_1_propagate_pipe_b <= mesh_6_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_2_io_in_control_0_shift_pipe_b <= mesh_7_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_2_io_in_control_0_dataflow_pipe_b <= mesh_7_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_2_io_in_control_0_propagate_pipe_b <= mesh_7_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_2_io_in_control_1_shift_pipe_b <= mesh_7_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_2_io_in_control_1_dataflow_pipe_b <= mesh_7_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_2_io_in_control_1_propagate_pipe_b <= mesh_7_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_2_io_in_control_0_shift_pipe_b <= mesh_8_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_2_io_in_control_0_dataflow_pipe_b <= mesh_8_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_2_io_in_control_0_propagate_pipe_b <= mesh_8_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_2_io_in_control_1_shift_pipe_b <= mesh_8_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_2_io_in_control_1_dataflow_pipe_b <= mesh_8_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_2_io_in_control_1_propagate_pipe_b <= mesh_8_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_2_io_in_control_0_shift_pipe_b <= mesh_9_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_2_io_in_control_0_dataflow_pipe_b <= mesh_9_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_2_io_in_control_0_propagate_pipe_b <= mesh_9_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_2_io_in_control_1_shift_pipe_b <= mesh_9_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_2_io_in_control_1_dataflow_pipe_b <= mesh_9_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_2_io_in_control_1_propagate_pipe_b <= mesh_9_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_2_io_in_control_0_shift_pipe_b <= mesh_10_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_2_io_in_control_0_dataflow_pipe_b <= mesh_10_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_2_io_in_control_0_propagate_pipe_b <= mesh_10_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_2_io_in_control_1_shift_pipe_b <= mesh_10_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_2_io_in_control_1_dataflow_pipe_b <= mesh_10_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_2_io_in_control_1_propagate_pipe_b <= mesh_10_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_2_io_in_control_0_shift_pipe_b <= mesh_11_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_2_io_in_control_0_dataflow_pipe_b <= mesh_11_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_2_io_in_control_0_propagate_pipe_b <= mesh_11_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_2_io_in_control_1_shift_pipe_b <= mesh_11_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_2_io_in_control_1_dataflow_pipe_b <= mesh_11_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_2_io_in_control_1_propagate_pipe_b <= mesh_11_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_2_io_in_control_0_shift_pipe_b <= mesh_12_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_2_io_in_control_0_dataflow_pipe_b <= mesh_12_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_2_io_in_control_0_propagate_pipe_b <= mesh_12_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_2_io_in_control_1_shift_pipe_b <= mesh_12_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_2_io_in_control_1_dataflow_pipe_b <= mesh_12_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_2_io_in_control_1_propagate_pipe_b <= mesh_12_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_2_io_in_control_0_shift_pipe_b <= mesh_13_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_2_io_in_control_0_dataflow_pipe_b <= mesh_13_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_2_io_in_control_0_propagate_pipe_b <= mesh_13_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_2_io_in_control_1_shift_pipe_b <= mesh_13_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_2_io_in_control_1_dataflow_pipe_b <= mesh_13_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_2_io_in_control_1_propagate_pipe_b <= mesh_13_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_2_io_in_control_0_shift_pipe_b <= mesh_14_2_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_2_io_in_control_0_dataflow_pipe_b <= mesh_14_2_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_2_io_in_control_0_propagate_pipe_b <= mesh_14_2_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_2_io_in_control_1_shift_pipe_b <= mesh_14_2_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_2_io_in_control_1_dataflow_pipe_b <= mesh_14_2_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_2_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_2_io_in_control_1_propagate_pipe_b <= mesh_14_2_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_3_io_in_control_0_shift_pipe_b <= io_in_control_3_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_3_io_in_control_0_dataflow_pipe_b <= io_in_control_3_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_3_io_in_control_0_propagate_pipe_b <= io_in_control_3_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_3_io_in_control_1_shift_pipe_b <= io_in_control_3_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_3_io_in_control_1_dataflow_pipe_b <= io_in_control_3_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_3_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_3_io_in_control_1_propagate_pipe_b <= io_in_control_3_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_3_io_in_control_0_shift_pipe_b <= mesh_0_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_3_io_in_control_0_dataflow_pipe_b <= mesh_0_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_3_io_in_control_0_propagate_pipe_b <= mesh_0_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_3_io_in_control_1_shift_pipe_b <= mesh_0_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_3_io_in_control_1_dataflow_pipe_b <= mesh_0_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_3_io_in_control_1_propagate_pipe_b <= mesh_0_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_3_io_in_control_0_shift_pipe_b <= mesh_1_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_3_io_in_control_0_dataflow_pipe_b <= mesh_1_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_3_io_in_control_0_propagate_pipe_b <= mesh_1_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_3_io_in_control_1_shift_pipe_b <= mesh_1_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_3_io_in_control_1_dataflow_pipe_b <= mesh_1_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_3_io_in_control_1_propagate_pipe_b <= mesh_1_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_3_io_in_control_0_shift_pipe_b <= mesh_2_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_3_io_in_control_0_dataflow_pipe_b <= mesh_2_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_3_io_in_control_0_propagate_pipe_b <= mesh_2_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_3_io_in_control_1_shift_pipe_b <= mesh_2_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_3_io_in_control_1_dataflow_pipe_b <= mesh_2_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_3_io_in_control_1_propagate_pipe_b <= mesh_2_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_3_io_in_control_0_shift_pipe_b <= mesh_3_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_3_io_in_control_0_dataflow_pipe_b <= mesh_3_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_3_io_in_control_0_propagate_pipe_b <= mesh_3_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_3_io_in_control_1_shift_pipe_b <= mesh_3_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_3_io_in_control_1_dataflow_pipe_b <= mesh_3_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_3_io_in_control_1_propagate_pipe_b <= mesh_3_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_3_io_in_control_0_shift_pipe_b <= mesh_4_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_3_io_in_control_0_dataflow_pipe_b <= mesh_4_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_3_io_in_control_0_propagate_pipe_b <= mesh_4_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_3_io_in_control_1_shift_pipe_b <= mesh_4_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_3_io_in_control_1_dataflow_pipe_b <= mesh_4_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_3_io_in_control_1_propagate_pipe_b <= mesh_4_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_3_io_in_control_0_shift_pipe_b <= mesh_5_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_3_io_in_control_0_dataflow_pipe_b <= mesh_5_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_3_io_in_control_0_propagate_pipe_b <= mesh_5_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_3_io_in_control_1_shift_pipe_b <= mesh_5_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_3_io_in_control_1_dataflow_pipe_b <= mesh_5_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_3_io_in_control_1_propagate_pipe_b <= mesh_5_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_3_io_in_control_0_shift_pipe_b <= mesh_6_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_3_io_in_control_0_dataflow_pipe_b <= mesh_6_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_3_io_in_control_0_propagate_pipe_b <= mesh_6_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_3_io_in_control_1_shift_pipe_b <= mesh_6_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_3_io_in_control_1_dataflow_pipe_b <= mesh_6_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_3_io_in_control_1_propagate_pipe_b <= mesh_6_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_3_io_in_control_0_shift_pipe_b <= mesh_7_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_3_io_in_control_0_dataflow_pipe_b <= mesh_7_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_3_io_in_control_0_propagate_pipe_b <= mesh_7_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_3_io_in_control_1_shift_pipe_b <= mesh_7_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_3_io_in_control_1_dataflow_pipe_b <= mesh_7_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_3_io_in_control_1_propagate_pipe_b <= mesh_7_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_3_io_in_control_0_shift_pipe_b <= mesh_8_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_3_io_in_control_0_dataflow_pipe_b <= mesh_8_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_3_io_in_control_0_propagate_pipe_b <= mesh_8_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_3_io_in_control_1_shift_pipe_b <= mesh_8_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_3_io_in_control_1_dataflow_pipe_b <= mesh_8_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_3_io_in_control_1_propagate_pipe_b <= mesh_8_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_3_io_in_control_0_shift_pipe_b <= mesh_9_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_3_io_in_control_0_dataflow_pipe_b <= mesh_9_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_3_io_in_control_0_propagate_pipe_b <= mesh_9_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_3_io_in_control_1_shift_pipe_b <= mesh_9_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_3_io_in_control_1_dataflow_pipe_b <= mesh_9_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_3_io_in_control_1_propagate_pipe_b <= mesh_9_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_3_io_in_control_0_shift_pipe_b <= mesh_10_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_3_io_in_control_0_dataflow_pipe_b <= mesh_10_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_3_io_in_control_0_propagate_pipe_b <= mesh_10_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_3_io_in_control_1_shift_pipe_b <= mesh_10_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_3_io_in_control_1_dataflow_pipe_b <= mesh_10_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_3_io_in_control_1_propagate_pipe_b <= mesh_10_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_3_io_in_control_0_shift_pipe_b <= mesh_11_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_3_io_in_control_0_dataflow_pipe_b <= mesh_11_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_3_io_in_control_0_propagate_pipe_b <= mesh_11_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_3_io_in_control_1_shift_pipe_b <= mesh_11_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_3_io_in_control_1_dataflow_pipe_b <= mesh_11_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_3_io_in_control_1_propagate_pipe_b <= mesh_11_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_3_io_in_control_0_shift_pipe_b <= mesh_12_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_3_io_in_control_0_dataflow_pipe_b <= mesh_12_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_3_io_in_control_0_propagate_pipe_b <= mesh_12_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_3_io_in_control_1_shift_pipe_b <= mesh_12_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_3_io_in_control_1_dataflow_pipe_b <= mesh_12_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_3_io_in_control_1_propagate_pipe_b <= mesh_12_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_3_io_in_control_0_shift_pipe_b <= mesh_13_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_3_io_in_control_0_dataflow_pipe_b <= mesh_13_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_3_io_in_control_0_propagate_pipe_b <= mesh_13_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_3_io_in_control_1_shift_pipe_b <= mesh_13_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_3_io_in_control_1_dataflow_pipe_b <= mesh_13_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_3_io_in_control_1_propagate_pipe_b <= mesh_13_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_3_io_in_control_0_shift_pipe_b <= mesh_14_3_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_3_io_in_control_0_dataflow_pipe_b <= mesh_14_3_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_3_io_in_control_0_propagate_pipe_b <= mesh_14_3_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_3_io_in_control_1_shift_pipe_b <= mesh_14_3_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_3_io_in_control_1_dataflow_pipe_b <= mesh_14_3_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_3_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_3_io_in_control_1_propagate_pipe_b <= mesh_14_3_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_4_io_in_control_0_shift_pipe_b <= io_in_control_4_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_4_io_in_control_0_dataflow_pipe_b <= io_in_control_4_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_4_io_in_control_0_propagate_pipe_b <= io_in_control_4_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_4_io_in_control_1_shift_pipe_b <= io_in_control_4_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_4_io_in_control_1_dataflow_pipe_b <= io_in_control_4_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_4_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_4_io_in_control_1_propagate_pipe_b <= io_in_control_4_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_4_io_in_control_0_shift_pipe_b <= mesh_0_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_4_io_in_control_0_dataflow_pipe_b <= mesh_0_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_4_io_in_control_0_propagate_pipe_b <= mesh_0_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_4_io_in_control_1_shift_pipe_b <= mesh_0_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_4_io_in_control_1_dataflow_pipe_b <= mesh_0_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_4_io_in_control_1_propagate_pipe_b <= mesh_0_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_4_io_in_control_0_shift_pipe_b <= mesh_1_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_4_io_in_control_0_dataflow_pipe_b <= mesh_1_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_4_io_in_control_0_propagate_pipe_b <= mesh_1_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_4_io_in_control_1_shift_pipe_b <= mesh_1_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_4_io_in_control_1_dataflow_pipe_b <= mesh_1_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_4_io_in_control_1_propagate_pipe_b <= mesh_1_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_4_io_in_control_0_shift_pipe_b <= mesh_2_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_4_io_in_control_0_dataflow_pipe_b <= mesh_2_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_4_io_in_control_0_propagate_pipe_b <= mesh_2_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_4_io_in_control_1_shift_pipe_b <= mesh_2_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_4_io_in_control_1_dataflow_pipe_b <= mesh_2_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_4_io_in_control_1_propagate_pipe_b <= mesh_2_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_4_io_in_control_0_shift_pipe_b <= mesh_3_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_4_io_in_control_0_dataflow_pipe_b <= mesh_3_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_4_io_in_control_0_propagate_pipe_b <= mesh_3_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_4_io_in_control_1_shift_pipe_b <= mesh_3_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_4_io_in_control_1_dataflow_pipe_b <= mesh_3_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_4_io_in_control_1_propagate_pipe_b <= mesh_3_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_4_io_in_control_0_shift_pipe_b <= mesh_4_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_4_io_in_control_0_dataflow_pipe_b <= mesh_4_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_4_io_in_control_0_propagate_pipe_b <= mesh_4_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_4_io_in_control_1_shift_pipe_b <= mesh_4_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_4_io_in_control_1_dataflow_pipe_b <= mesh_4_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_4_io_in_control_1_propagate_pipe_b <= mesh_4_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_4_io_in_control_0_shift_pipe_b <= mesh_5_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_4_io_in_control_0_dataflow_pipe_b <= mesh_5_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_4_io_in_control_0_propagate_pipe_b <= mesh_5_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_4_io_in_control_1_shift_pipe_b <= mesh_5_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_4_io_in_control_1_dataflow_pipe_b <= mesh_5_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_4_io_in_control_1_propagate_pipe_b <= mesh_5_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_4_io_in_control_0_shift_pipe_b <= mesh_6_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_4_io_in_control_0_dataflow_pipe_b <= mesh_6_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_4_io_in_control_0_propagate_pipe_b <= mesh_6_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_4_io_in_control_1_shift_pipe_b <= mesh_6_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_4_io_in_control_1_dataflow_pipe_b <= mesh_6_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_4_io_in_control_1_propagate_pipe_b <= mesh_6_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_4_io_in_control_0_shift_pipe_b <= mesh_7_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_4_io_in_control_0_dataflow_pipe_b <= mesh_7_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_4_io_in_control_0_propagate_pipe_b <= mesh_7_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_4_io_in_control_1_shift_pipe_b <= mesh_7_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_4_io_in_control_1_dataflow_pipe_b <= mesh_7_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_4_io_in_control_1_propagate_pipe_b <= mesh_7_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_4_io_in_control_0_shift_pipe_b <= mesh_8_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_4_io_in_control_0_dataflow_pipe_b <= mesh_8_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_4_io_in_control_0_propagate_pipe_b <= mesh_8_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_4_io_in_control_1_shift_pipe_b <= mesh_8_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_4_io_in_control_1_dataflow_pipe_b <= mesh_8_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_4_io_in_control_1_propagate_pipe_b <= mesh_8_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_4_io_in_control_0_shift_pipe_b <= mesh_9_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_4_io_in_control_0_dataflow_pipe_b <= mesh_9_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_4_io_in_control_0_propagate_pipe_b <= mesh_9_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_4_io_in_control_1_shift_pipe_b <= mesh_9_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_4_io_in_control_1_dataflow_pipe_b <= mesh_9_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_4_io_in_control_1_propagate_pipe_b <= mesh_9_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_4_io_in_control_0_shift_pipe_b <= mesh_10_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_4_io_in_control_0_dataflow_pipe_b <= mesh_10_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_4_io_in_control_0_propagate_pipe_b <= mesh_10_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_4_io_in_control_1_shift_pipe_b <= mesh_10_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_4_io_in_control_1_dataflow_pipe_b <= mesh_10_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_4_io_in_control_1_propagate_pipe_b <= mesh_10_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_4_io_in_control_0_shift_pipe_b <= mesh_11_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_4_io_in_control_0_dataflow_pipe_b <= mesh_11_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_4_io_in_control_0_propagate_pipe_b <= mesh_11_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_4_io_in_control_1_shift_pipe_b <= mesh_11_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_4_io_in_control_1_dataflow_pipe_b <= mesh_11_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_4_io_in_control_1_propagate_pipe_b <= mesh_11_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_4_io_in_control_0_shift_pipe_b <= mesh_12_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_4_io_in_control_0_dataflow_pipe_b <= mesh_12_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_4_io_in_control_0_propagate_pipe_b <= mesh_12_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_4_io_in_control_1_shift_pipe_b <= mesh_12_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_4_io_in_control_1_dataflow_pipe_b <= mesh_12_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_4_io_in_control_1_propagate_pipe_b <= mesh_12_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_4_io_in_control_0_shift_pipe_b <= mesh_13_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_4_io_in_control_0_dataflow_pipe_b <= mesh_13_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_4_io_in_control_0_propagate_pipe_b <= mesh_13_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_4_io_in_control_1_shift_pipe_b <= mesh_13_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_4_io_in_control_1_dataflow_pipe_b <= mesh_13_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_4_io_in_control_1_propagate_pipe_b <= mesh_13_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_4_io_in_control_0_shift_pipe_b <= mesh_14_4_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_4_io_in_control_0_dataflow_pipe_b <= mesh_14_4_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_4_io_in_control_0_propagate_pipe_b <= mesh_14_4_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_4_io_in_control_1_shift_pipe_b <= mesh_14_4_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_4_io_in_control_1_dataflow_pipe_b <= mesh_14_4_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_4_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_4_io_in_control_1_propagate_pipe_b <= mesh_14_4_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_5_io_in_control_0_shift_pipe_b <= io_in_control_5_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_5_io_in_control_0_dataflow_pipe_b <= io_in_control_5_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_5_io_in_control_0_propagate_pipe_b <= io_in_control_5_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_5_io_in_control_1_shift_pipe_b <= io_in_control_5_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_5_io_in_control_1_dataflow_pipe_b <= io_in_control_5_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_5_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_5_io_in_control_1_propagate_pipe_b <= io_in_control_5_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_5_io_in_control_0_shift_pipe_b <= mesh_0_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_5_io_in_control_0_dataflow_pipe_b <= mesh_0_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_5_io_in_control_0_propagate_pipe_b <= mesh_0_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_5_io_in_control_1_shift_pipe_b <= mesh_0_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_5_io_in_control_1_dataflow_pipe_b <= mesh_0_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_5_io_in_control_1_propagate_pipe_b <= mesh_0_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_5_io_in_control_0_shift_pipe_b <= mesh_1_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_5_io_in_control_0_dataflow_pipe_b <= mesh_1_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_5_io_in_control_0_propagate_pipe_b <= mesh_1_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_5_io_in_control_1_shift_pipe_b <= mesh_1_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_5_io_in_control_1_dataflow_pipe_b <= mesh_1_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_5_io_in_control_1_propagate_pipe_b <= mesh_1_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_5_io_in_control_0_shift_pipe_b <= mesh_2_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_5_io_in_control_0_dataflow_pipe_b <= mesh_2_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_5_io_in_control_0_propagate_pipe_b <= mesh_2_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_5_io_in_control_1_shift_pipe_b <= mesh_2_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_5_io_in_control_1_dataflow_pipe_b <= mesh_2_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_5_io_in_control_1_propagate_pipe_b <= mesh_2_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_5_io_in_control_0_shift_pipe_b <= mesh_3_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_5_io_in_control_0_dataflow_pipe_b <= mesh_3_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_5_io_in_control_0_propagate_pipe_b <= mesh_3_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_5_io_in_control_1_shift_pipe_b <= mesh_3_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_5_io_in_control_1_dataflow_pipe_b <= mesh_3_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_5_io_in_control_1_propagate_pipe_b <= mesh_3_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_5_io_in_control_0_shift_pipe_b <= mesh_4_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_5_io_in_control_0_dataflow_pipe_b <= mesh_4_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_5_io_in_control_0_propagate_pipe_b <= mesh_4_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_5_io_in_control_1_shift_pipe_b <= mesh_4_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_5_io_in_control_1_dataflow_pipe_b <= mesh_4_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_5_io_in_control_1_propagate_pipe_b <= mesh_4_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_5_io_in_control_0_shift_pipe_b <= mesh_5_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_5_io_in_control_0_dataflow_pipe_b <= mesh_5_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_5_io_in_control_0_propagate_pipe_b <= mesh_5_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_5_io_in_control_1_shift_pipe_b <= mesh_5_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_5_io_in_control_1_dataflow_pipe_b <= mesh_5_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_5_io_in_control_1_propagate_pipe_b <= mesh_5_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_5_io_in_control_0_shift_pipe_b <= mesh_6_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_5_io_in_control_0_dataflow_pipe_b <= mesh_6_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_5_io_in_control_0_propagate_pipe_b <= mesh_6_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_5_io_in_control_1_shift_pipe_b <= mesh_6_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_5_io_in_control_1_dataflow_pipe_b <= mesh_6_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_5_io_in_control_1_propagate_pipe_b <= mesh_6_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_5_io_in_control_0_shift_pipe_b <= mesh_7_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_5_io_in_control_0_dataflow_pipe_b <= mesh_7_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_5_io_in_control_0_propagate_pipe_b <= mesh_7_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_5_io_in_control_1_shift_pipe_b <= mesh_7_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_5_io_in_control_1_dataflow_pipe_b <= mesh_7_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_5_io_in_control_1_propagate_pipe_b <= mesh_7_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_5_io_in_control_0_shift_pipe_b <= mesh_8_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_5_io_in_control_0_dataflow_pipe_b <= mesh_8_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_5_io_in_control_0_propagate_pipe_b <= mesh_8_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_5_io_in_control_1_shift_pipe_b <= mesh_8_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_5_io_in_control_1_dataflow_pipe_b <= mesh_8_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_5_io_in_control_1_propagate_pipe_b <= mesh_8_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_5_io_in_control_0_shift_pipe_b <= mesh_9_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_5_io_in_control_0_dataflow_pipe_b <= mesh_9_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_5_io_in_control_0_propagate_pipe_b <= mesh_9_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_5_io_in_control_1_shift_pipe_b <= mesh_9_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_5_io_in_control_1_dataflow_pipe_b <= mesh_9_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_5_io_in_control_1_propagate_pipe_b <= mesh_9_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_5_io_in_control_0_shift_pipe_b <= mesh_10_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_5_io_in_control_0_dataflow_pipe_b <= mesh_10_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_5_io_in_control_0_propagate_pipe_b <= mesh_10_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_5_io_in_control_1_shift_pipe_b <= mesh_10_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_5_io_in_control_1_dataflow_pipe_b <= mesh_10_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_5_io_in_control_1_propagate_pipe_b <= mesh_10_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_5_io_in_control_0_shift_pipe_b <= mesh_11_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_5_io_in_control_0_dataflow_pipe_b <= mesh_11_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_5_io_in_control_0_propagate_pipe_b <= mesh_11_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_5_io_in_control_1_shift_pipe_b <= mesh_11_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_5_io_in_control_1_dataflow_pipe_b <= mesh_11_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_5_io_in_control_1_propagate_pipe_b <= mesh_11_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_5_io_in_control_0_shift_pipe_b <= mesh_12_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_5_io_in_control_0_dataflow_pipe_b <= mesh_12_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_5_io_in_control_0_propagate_pipe_b <= mesh_12_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_5_io_in_control_1_shift_pipe_b <= mesh_12_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_5_io_in_control_1_dataflow_pipe_b <= mesh_12_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_5_io_in_control_1_propagate_pipe_b <= mesh_12_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_5_io_in_control_0_shift_pipe_b <= mesh_13_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_5_io_in_control_0_dataflow_pipe_b <= mesh_13_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_5_io_in_control_0_propagate_pipe_b <= mesh_13_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_5_io_in_control_1_shift_pipe_b <= mesh_13_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_5_io_in_control_1_dataflow_pipe_b <= mesh_13_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_5_io_in_control_1_propagate_pipe_b <= mesh_13_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_5_io_in_control_0_shift_pipe_b <= mesh_14_5_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_5_io_in_control_0_dataflow_pipe_b <= mesh_14_5_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_5_io_in_control_0_propagate_pipe_b <= mesh_14_5_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_5_io_in_control_1_shift_pipe_b <= mesh_14_5_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_5_io_in_control_1_dataflow_pipe_b <= mesh_14_5_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_5_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_5_io_in_control_1_propagate_pipe_b <= mesh_14_5_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_6_io_in_control_0_shift_pipe_b <= io_in_control_6_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_6_io_in_control_0_dataflow_pipe_b <= io_in_control_6_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_6_io_in_control_0_propagate_pipe_b <= io_in_control_6_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_6_io_in_control_1_shift_pipe_b <= io_in_control_6_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_6_io_in_control_1_dataflow_pipe_b <= io_in_control_6_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_6_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_6_io_in_control_1_propagate_pipe_b <= io_in_control_6_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_6_io_in_control_0_shift_pipe_b <= mesh_0_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_6_io_in_control_0_dataflow_pipe_b <= mesh_0_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_6_io_in_control_0_propagate_pipe_b <= mesh_0_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_6_io_in_control_1_shift_pipe_b <= mesh_0_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_6_io_in_control_1_dataflow_pipe_b <= mesh_0_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_6_io_in_control_1_propagate_pipe_b <= mesh_0_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_6_io_in_control_0_shift_pipe_b <= mesh_1_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_6_io_in_control_0_dataflow_pipe_b <= mesh_1_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_6_io_in_control_0_propagate_pipe_b <= mesh_1_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_6_io_in_control_1_shift_pipe_b <= mesh_1_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_6_io_in_control_1_dataflow_pipe_b <= mesh_1_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_6_io_in_control_1_propagate_pipe_b <= mesh_1_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_6_io_in_control_0_shift_pipe_b <= mesh_2_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_6_io_in_control_0_dataflow_pipe_b <= mesh_2_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_6_io_in_control_0_propagate_pipe_b <= mesh_2_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_6_io_in_control_1_shift_pipe_b <= mesh_2_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_6_io_in_control_1_dataflow_pipe_b <= mesh_2_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_6_io_in_control_1_propagate_pipe_b <= mesh_2_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_6_io_in_control_0_shift_pipe_b <= mesh_3_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_6_io_in_control_0_dataflow_pipe_b <= mesh_3_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_6_io_in_control_0_propagate_pipe_b <= mesh_3_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_6_io_in_control_1_shift_pipe_b <= mesh_3_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_6_io_in_control_1_dataflow_pipe_b <= mesh_3_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_6_io_in_control_1_propagate_pipe_b <= mesh_3_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_6_io_in_control_0_shift_pipe_b <= mesh_4_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_6_io_in_control_0_dataflow_pipe_b <= mesh_4_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_6_io_in_control_0_propagate_pipe_b <= mesh_4_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_6_io_in_control_1_shift_pipe_b <= mesh_4_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_6_io_in_control_1_dataflow_pipe_b <= mesh_4_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_6_io_in_control_1_propagate_pipe_b <= mesh_4_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_6_io_in_control_0_shift_pipe_b <= mesh_5_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_6_io_in_control_0_dataflow_pipe_b <= mesh_5_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_6_io_in_control_0_propagate_pipe_b <= mesh_5_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_6_io_in_control_1_shift_pipe_b <= mesh_5_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_6_io_in_control_1_dataflow_pipe_b <= mesh_5_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_6_io_in_control_1_propagate_pipe_b <= mesh_5_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_6_io_in_control_0_shift_pipe_b <= mesh_6_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_6_io_in_control_0_dataflow_pipe_b <= mesh_6_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_6_io_in_control_0_propagate_pipe_b <= mesh_6_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_6_io_in_control_1_shift_pipe_b <= mesh_6_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_6_io_in_control_1_dataflow_pipe_b <= mesh_6_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_6_io_in_control_1_propagate_pipe_b <= mesh_6_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_6_io_in_control_0_shift_pipe_b <= mesh_7_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_6_io_in_control_0_dataflow_pipe_b <= mesh_7_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_6_io_in_control_0_propagate_pipe_b <= mesh_7_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_6_io_in_control_1_shift_pipe_b <= mesh_7_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_6_io_in_control_1_dataflow_pipe_b <= mesh_7_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_6_io_in_control_1_propagate_pipe_b <= mesh_7_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_6_io_in_control_0_shift_pipe_b <= mesh_8_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_6_io_in_control_0_dataflow_pipe_b <= mesh_8_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_6_io_in_control_0_propagate_pipe_b <= mesh_8_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_6_io_in_control_1_shift_pipe_b <= mesh_8_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_6_io_in_control_1_dataflow_pipe_b <= mesh_8_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_6_io_in_control_1_propagate_pipe_b <= mesh_8_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_6_io_in_control_0_shift_pipe_b <= mesh_9_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_6_io_in_control_0_dataflow_pipe_b <= mesh_9_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_6_io_in_control_0_propagate_pipe_b <= mesh_9_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_6_io_in_control_1_shift_pipe_b <= mesh_9_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_6_io_in_control_1_dataflow_pipe_b <= mesh_9_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_6_io_in_control_1_propagate_pipe_b <= mesh_9_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_6_io_in_control_0_shift_pipe_b <= mesh_10_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_6_io_in_control_0_dataflow_pipe_b <= mesh_10_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_6_io_in_control_0_propagate_pipe_b <= mesh_10_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_6_io_in_control_1_shift_pipe_b <= mesh_10_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_6_io_in_control_1_dataflow_pipe_b <= mesh_10_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_6_io_in_control_1_propagate_pipe_b <= mesh_10_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_6_io_in_control_0_shift_pipe_b <= mesh_11_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_6_io_in_control_0_dataflow_pipe_b <= mesh_11_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_6_io_in_control_0_propagate_pipe_b <= mesh_11_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_6_io_in_control_1_shift_pipe_b <= mesh_11_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_6_io_in_control_1_dataflow_pipe_b <= mesh_11_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_6_io_in_control_1_propagate_pipe_b <= mesh_11_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_6_io_in_control_0_shift_pipe_b <= mesh_12_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_6_io_in_control_0_dataflow_pipe_b <= mesh_12_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_6_io_in_control_0_propagate_pipe_b <= mesh_12_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_6_io_in_control_1_shift_pipe_b <= mesh_12_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_6_io_in_control_1_dataflow_pipe_b <= mesh_12_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_6_io_in_control_1_propagate_pipe_b <= mesh_12_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_6_io_in_control_0_shift_pipe_b <= mesh_13_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_6_io_in_control_0_dataflow_pipe_b <= mesh_13_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_6_io_in_control_0_propagate_pipe_b <= mesh_13_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_6_io_in_control_1_shift_pipe_b <= mesh_13_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_6_io_in_control_1_dataflow_pipe_b <= mesh_13_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_6_io_in_control_1_propagate_pipe_b <= mesh_13_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_6_io_in_control_0_shift_pipe_b <= mesh_14_6_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_6_io_in_control_0_dataflow_pipe_b <= mesh_14_6_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_6_io_in_control_0_propagate_pipe_b <= mesh_14_6_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_6_io_in_control_1_shift_pipe_b <= mesh_14_6_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_6_io_in_control_1_dataflow_pipe_b <= mesh_14_6_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_6_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_6_io_in_control_1_propagate_pipe_b <= mesh_14_6_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_7_io_in_control_0_shift_pipe_b <= io_in_control_7_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_7_io_in_control_0_dataflow_pipe_b <= io_in_control_7_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_7_io_in_control_0_propagate_pipe_b <= io_in_control_7_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_7_io_in_control_1_shift_pipe_b <= io_in_control_7_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_7_io_in_control_1_dataflow_pipe_b <= io_in_control_7_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_7_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_7_io_in_control_1_propagate_pipe_b <= io_in_control_7_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_7_io_in_control_0_shift_pipe_b <= mesh_0_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_7_io_in_control_0_dataflow_pipe_b <= mesh_0_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_7_io_in_control_0_propagate_pipe_b <= mesh_0_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_7_io_in_control_1_shift_pipe_b <= mesh_0_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_7_io_in_control_1_dataflow_pipe_b <= mesh_0_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_7_io_in_control_1_propagate_pipe_b <= mesh_0_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_7_io_in_control_0_shift_pipe_b <= mesh_1_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_7_io_in_control_0_dataflow_pipe_b <= mesh_1_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_7_io_in_control_0_propagate_pipe_b <= mesh_1_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_7_io_in_control_1_shift_pipe_b <= mesh_1_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_7_io_in_control_1_dataflow_pipe_b <= mesh_1_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_7_io_in_control_1_propagate_pipe_b <= mesh_1_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_7_io_in_control_0_shift_pipe_b <= mesh_2_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_7_io_in_control_0_dataflow_pipe_b <= mesh_2_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_7_io_in_control_0_propagate_pipe_b <= mesh_2_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_7_io_in_control_1_shift_pipe_b <= mesh_2_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_7_io_in_control_1_dataflow_pipe_b <= mesh_2_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_7_io_in_control_1_propagate_pipe_b <= mesh_2_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_7_io_in_control_0_shift_pipe_b <= mesh_3_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_7_io_in_control_0_dataflow_pipe_b <= mesh_3_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_7_io_in_control_0_propagate_pipe_b <= mesh_3_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_7_io_in_control_1_shift_pipe_b <= mesh_3_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_7_io_in_control_1_dataflow_pipe_b <= mesh_3_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_7_io_in_control_1_propagate_pipe_b <= mesh_3_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_7_io_in_control_0_shift_pipe_b <= mesh_4_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_7_io_in_control_0_dataflow_pipe_b <= mesh_4_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_7_io_in_control_0_propagate_pipe_b <= mesh_4_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_7_io_in_control_1_shift_pipe_b <= mesh_4_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_7_io_in_control_1_dataflow_pipe_b <= mesh_4_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_7_io_in_control_1_propagate_pipe_b <= mesh_4_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_7_io_in_control_0_shift_pipe_b <= mesh_5_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_7_io_in_control_0_dataflow_pipe_b <= mesh_5_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_7_io_in_control_0_propagate_pipe_b <= mesh_5_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_7_io_in_control_1_shift_pipe_b <= mesh_5_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_7_io_in_control_1_dataflow_pipe_b <= mesh_5_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_7_io_in_control_1_propagate_pipe_b <= mesh_5_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_7_io_in_control_0_shift_pipe_b <= mesh_6_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_7_io_in_control_0_dataflow_pipe_b <= mesh_6_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_7_io_in_control_0_propagate_pipe_b <= mesh_6_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_7_io_in_control_1_shift_pipe_b <= mesh_6_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_7_io_in_control_1_dataflow_pipe_b <= mesh_6_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_7_io_in_control_1_propagate_pipe_b <= mesh_6_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_7_io_in_control_0_shift_pipe_b <= mesh_7_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_7_io_in_control_0_dataflow_pipe_b <= mesh_7_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_7_io_in_control_0_propagate_pipe_b <= mesh_7_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_7_io_in_control_1_shift_pipe_b <= mesh_7_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_7_io_in_control_1_dataflow_pipe_b <= mesh_7_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_7_io_in_control_1_propagate_pipe_b <= mesh_7_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_7_io_in_control_0_shift_pipe_b <= mesh_8_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_7_io_in_control_0_dataflow_pipe_b <= mesh_8_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_7_io_in_control_0_propagate_pipe_b <= mesh_8_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_7_io_in_control_1_shift_pipe_b <= mesh_8_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_7_io_in_control_1_dataflow_pipe_b <= mesh_8_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_7_io_in_control_1_propagate_pipe_b <= mesh_8_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_7_io_in_control_0_shift_pipe_b <= mesh_9_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_7_io_in_control_0_dataflow_pipe_b <= mesh_9_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_7_io_in_control_0_propagate_pipe_b <= mesh_9_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_7_io_in_control_1_shift_pipe_b <= mesh_9_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_7_io_in_control_1_dataflow_pipe_b <= mesh_9_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_7_io_in_control_1_propagate_pipe_b <= mesh_9_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_7_io_in_control_0_shift_pipe_b <= mesh_10_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_7_io_in_control_0_dataflow_pipe_b <= mesh_10_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_7_io_in_control_0_propagate_pipe_b <= mesh_10_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_7_io_in_control_1_shift_pipe_b <= mesh_10_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_7_io_in_control_1_dataflow_pipe_b <= mesh_10_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_7_io_in_control_1_propagate_pipe_b <= mesh_10_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_7_io_in_control_0_shift_pipe_b <= mesh_11_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_7_io_in_control_0_dataflow_pipe_b <= mesh_11_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_7_io_in_control_0_propagate_pipe_b <= mesh_11_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_7_io_in_control_1_shift_pipe_b <= mesh_11_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_7_io_in_control_1_dataflow_pipe_b <= mesh_11_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_7_io_in_control_1_propagate_pipe_b <= mesh_11_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_7_io_in_control_0_shift_pipe_b <= mesh_12_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_7_io_in_control_0_dataflow_pipe_b <= mesh_12_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_7_io_in_control_0_propagate_pipe_b <= mesh_12_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_7_io_in_control_1_shift_pipe_b <= mesh_12_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_7_io_in_control_1_dataflow_pipe_b <= mesh_12_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_7_io_in_control_1_propagate_pipe_b <= mesh_12_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_7_io_in_control_0_shift_pipe_b <= mesh_13_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_7_io_in_control_0_dataflow_pipe_b <= mesh_13_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_7_io_in_control_0_propagate_pipe_b <= mesh_13_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_7_io_in_control_1_shift_pipe_b <= mesh_13_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_7_io_in_control_1_dataflow_pipe_b <= mesh_13_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_7_io_in_control_1_propagate_pipe_b <= mesh_13_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_7_io_in_control_0_shift_pipe_b <= mesh_14_7_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_7_io_in_control_0_dataflow_pipe_b <= mesh_14_7_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_7_io_in_control_0_propagate_pipe_b <= mesh_14_7_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_7_io_in_control_1_shift_pipe_b <= mesh_14_7_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_7_io_in_control_1_dataflow_pipe_b <= mesh_14_7_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_7_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_7_io_in_control_1_propagate_pipe_b <= mesh_14_7_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_8_io_in_control_0_shift_pipe_b <= io_in_control_8_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_8_io_in_control_0_dataflow_pipe_b <= io_in_control_8_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_8_io_in_control_0_propagate_pipe_b <= io_in_control_8_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_8_io_in_control_1_shift_pipe_b <= io_in_control_8_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_8_io_in_control_1_dataflow_pipe_b <= io_in_control_8_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_8_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_8_io_in_control_1_propagate_pipe_b <= io_in_control_8_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_8_io_in_control_0_shift_pipe_b <= mesh_0_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_8_io_in_control_0_dataflow_pipe_b <= mesh_0_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_8_io_in_control_0_propagate_pipe_b <= mesh_0_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_8_io_in_control_1_shift_pipe_b <= mesh_0_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_8_io_in_control_1_dataflow_pipe_b <= mesh_0_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_8_io_in_control_1_propagate_pipe_b <= mesh_0_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_8_io_in_control_0_shift_pipe_b <= mesh_1_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_8_io_in_control_0_dataflow_pipe_b <= mesh_1_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_8_io_in_control_0_propagate_pipe_b <= mesh_1_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_8_io_in_control_1_shift_pipe_b <= mesh_1_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_8_io_in_control_1_dataflow_pipe_b <= mesh_1_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_8_io_in_control_1_propagate_pipe_b <= mesh_1_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_8_io_in_control_0_shift_pipe_b <= mesh_2_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_8_io_in_control_0_dataflow_pipe_b <= mesh_2_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_8_io_in_control_0_propagate_pipe_b <= mesh_2_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_8_io_in_control_1_shift_pipe_b <= mesh_2_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_8_io_in_control_1_dataflow_pipe_b <= mesh_2_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_8_io_in_control_1_propagate_pipe_b <= mesh_2_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_8_io_in_control_0_shift_pipe_b <= mesh_3_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_8_io_in_control_0_dataflow_pipe_b <= mesh_3_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_8_io_in_control_0_propagate_pipe_b <= mesh_3_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_8_io_in_control_1_shift_pipe_b <= mesh_3_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_8_io_in_control_1_dataflow_pipe_b <= mesh_3_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_8_io_in_control_1_propagate_pipe_b <= mesh_3_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_8_io_in_control_0_shift_pipe_b <= mesh_4_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_8_io_in_control_0_dataflow_pipe_b <= mesh_4_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_8_io_in_control_0_propagate_pipe_b <= mesh_4_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_8_io_in_control_1_shift_pipe_b <= mesh_4_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_8_io_in_control_1_dataflow_pipe_b <= mesh_4_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_8_io_in_control_1_propagate_pipe_b <= mesh_4_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_8_io_in_control_0_shift_pipe_b <= mesh_5_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_8_io_in_control_0_dataflow_pipe_b <= mesh_5_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_8_io_in_control_0_propagate_pipe_b <= mesh_5_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_8_io_in_control_1_shift_pipe_b <= mesh_5_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_8_io_in_control_1_dataflow_pipe_b <= mesh_5_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_8_io_in_control_1_propagate_pipe_b <= mesh_5_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_8_io_in_control_0_shift_pipe_b <= mesh_6_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_8_io_in_control_0_dataflow_pipe_b <= mesh_6_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_8_io_in_control_0_propagate_pipe_b <= mesh_6_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_8_io_in_control_1_shift_pipe_b <= mesh_6_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_8_io_in_control_1_dataflow_pipe_b <= mesh_6_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_8_io_in_control_1_propagate_pipe_b <= mesh_6_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_8_io_in_control_0_shift_pipe_b <= mesh_7_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_8_io_in_control_0_dataflow_pipe_b <= mesh_7_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_8_io_in_control_0_propagate_pipe_b <= mesh_7_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_8_io_in_control_1_shift_pipe_b <= mesh_7_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_8_io_in_control_1_dataflow_pipe_b <= mesh_7_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_8_io_in_control_1_propagate_pipe_b <= mesh_7_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_8_io_in_control_0_shift_pipe_b <= mesh_8_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_8_io_in_control_0_dataflow_pipe_b <= mesh_8_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_8_io_in_control_0_propagate_pipe_b <= mesh_8_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_8_io_in_control_1_shift_pipe_b <= mesh_8_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_8_io_in_control_1_dataflow_pipe_b <= mesh_8_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_8_io_in_control_1_propagate_pipe_b <= mesh_8_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_8_io_in_control_0_shift_pipe_b <= mesh_9_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_8_io_in_control_0_dataflow_pipe_b <= mesh_9_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_8_io_in_control_0_propagate_pipe_b <= mesh_9_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_8_io_in_control_1_shift_pipe_b <= mesh_9_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_8_io_in_control_1_dataflow_pipe_b <= mesh_9_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_8_io_in_control_1_propagate_pipe_b <= mesh_9_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_8_io_in_control_0_shift_pipe_b <= mesh_10_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_8_io_in_control_0_dataflow_pipe_b <= mesh_10_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_8_io_in_control_0_propagate_pipe_b <= mesh_10_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_8_io_in_control_1_shift_pipe_b <= mesh_10_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_8_io_in_control_1_dataflow_pipe_b <= mesh_10_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_8_io_in_control_1_propagate_pipe_b <= mesh_10_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_8_io_in_control_0_shift_pipe_b <= mesh_11_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_8_io_in_control_0_dataflow_pipe_b <= mesh_11_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_8_io_in_control_0_propagate_pipe_b <= mesh_11_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_8_io_in_control_1_shift_pipe_b <= mesh_11_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_8_io_in_control_1_dataflow_pipe_b <= mesh_11_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_8_io_in_control_1_propagate_pipe_b <= mesh_11_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_8_io_in_control_0_shift_pipe_b <= mesh_12_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_8_io_in_control_0_dataflow_pipe_b <= mesh_12_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_8_io_in_control_0_propagate_pipe_b <= mesh_12_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_8_io_in_control_1_shift_pipe_b <= mesh_12_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_8_io_in_control_1_dataflow_pipe_b <= mesh_12_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_8_io_in_control_1_propagate_pipe_b <= mesh_12_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_8_io_in_control_0_shift_pipe_b <= mesh_13_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_8_io_in_control_0_dataflow_pipe_b <= mesh_13_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_8_io_in_control_0_propagate_pipe_b <= mesh_13_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_8_io_in_control_1_shift_pipe_b <= mesh_13_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_8_io_in_control_1_dataflow_pipe_b <= mesh_13_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_8_io_in_control_1_propagate_pipe_b <= mesh_13_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_8_io_in_control_0_shift_pipe_b <= mesh_14_8_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_8_io_in_control_0_dataflow_pipe_b <= mesh_14_8_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_8_io_in_control_0_propagate_pipe_b <= mesh_14_8_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_8_io_in_control_1_shift_pipe_b <= mesh_14_8_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_8_io_in_control_1_dataflow_pipe_b <= mesh_14_8_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_8_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_8_io_in_control_1_propagate_pipe_b <= mesh_14_8_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_9_io_in_control_0_shift_pipe_b <= io_in_control_9_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_9_io_in_control_0_dataflow_pipe_b <= io_in_control_9_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_9_io_in_control_0_propagate_pipe_b <= io_in_control_9_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_9_io_in_control_1_shift_pipe_b <= io_in_control_9_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_9_io_in_control_1_dataflow_pipe_b <= io_in_control_9_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_9_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_9_io_in_control_1_propagate_pipe_b <= io_in_control_9_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_9_io_in_control_0_shift_pipe_b <= mesh_0_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_9_io_in_control_0_dataflow_pipe_b <= mesh_0_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_9_io_in_control_0_propagate_pipe_b <= mesh_0_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_9_io_in_control_1_shift_pipe_b <= mesh_0_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_9_io_in_control_1_dataflow_pipe_b <= mesh_0_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_9_io_in_control_1_propagate_pipe_b <= mesh_0_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_9_io_in_control_0_shift_pipe_b <= mesh_1_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_9_io_in_control_0_dataflow_pipe_b <= mesh_1_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_9_io_in_control_0_propagate_pipe_b <= mesh_1_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_9_io_in_control_1_shift_pipe_b <= mesh_1_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_9_io_in_control_1_dataflow_pipe_b <= mesh_1_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_9_io_in_control_1_propagate_pipe_b <= mesh_1_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_9_io_in_control_0_shift_pipe_b <= mesh_2_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_9_io_in_control_0_dataflow_pipe_b <= mesh_2_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_9_io_in_control_0_propagate_pipe_b <= mesh_2_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_9_io_in_control_1_shift_pipe_b <= mesh_2_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_9_io_in_control_1_dataflow_pipe_b <= mesh_2_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_9_io_in_control_1_propagate_pipe_b <= mesh_2_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_9_io_in_control_0_shift_pipe_b <= mesh_3_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_9_io_in_control_0_dataflow_pipe_b <= mesh_3_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_9_io_in_control_0_propagate_pipe_b <= mesh_3_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_9_io_in_control_1_shift_pipe_b <= mesh_3_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_9_io_in_control_1_dataflow_pipe_b <= mesh_3_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_9_io_in_control_1_propagate_pipe_b <= mesh_3_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_9_io_in_control_0_shift_pipe_b <= mesh_4_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_9_io_in_control_0_dataflow_pipe_b <= mesh_4_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_9_io_in_control_0_propagate_pipe_b <= mesh_4_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_9_io_in_control_1_shift_pipe_b <= mesh_4_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_9_io_in_control_1_dataflow_pipe_b <= mesh_4_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_9_io_in_control_1_propagate_pipe_b <= mesh_4_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_9_io_in_control_0_shift_pipe_b <= mesh_5_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_9_io_in_control_0_dataflow_pipe_b <= mesh_5_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_9_io_in_control_0_propagate_pipe_b <= mesh_5_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_9_io_in_control_1_shift_pipe_b <= mesh_5_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_9_io_in_control_1_dataflow_pipe_b <= mesh_5_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_9_io_in_control_1_propagate_pipe_b <= mesh_5_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_9_io_in_control_0_shift_pipe_b <= mesh_6_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_9_io_in_control_0_dataflow_pipe_b <= mesh_6_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_9_io_in_control_0_propagate_pipe_b <= mesh_6_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_9_io_in_control_1_shift_pipe_b <= mesh_6_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_9_io_in_control_1_dataflow_pipe_b <= mesh_6_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_9_io_in_control_1_propagate_pipe_b <= mesh_6_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_9_io_in_control_0_shift_pipe_b <= mesh_7_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_9_io_in_control_0_dataflow_pipe_b <= mesh_7_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_9_io_in_control_0_propagate_pipe_b <= mesh_7_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_9_io_in_control_1_shift_pipe_b <= mesh_7_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_9_io_in_control_1_dataflow_pipe_b <= mesh_7_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_9_io_in_control_1_propagate_pipe_b <= mesh_7_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_9_io_in_control_0_shift_pipe_b <= mesh_8_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_9_io_in_control_0_dataflow_pipe_b <= mesh_8_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_9_io_in_control_0_propagate_pipe_b <= mesh_8_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_9_io_in_control_1_shift_pipe_b <= mesh_8_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_9_io_in_control_1_dataflow_pipe_b <= mesh_8_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_9_io_in_control_1_propagate_pipe_b <= mesh_8_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_9_io_in_control_0_shift_pipe_b <= mesh_9_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_9_io_in_control_0_dataflow_pipe_b <= mesh_9_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_9_io_in_control_0_propagate_pipe_b <= mesh_9_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_9_io_in_control_1_shift_pipe_b <= mesh_9_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_9_io_in_control_1_dataflow_pipe_b <= mesh_9_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_9_io_in_control_1_propagate_pipe_b <= mesh_9_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_9_io_in_control_0_shift_pipe_b <= mesh_10_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_9_io_in_control_0_dataflow_pipe_b <= mesh_10_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_9_io_in_control_0_propagate_pipe_b <= mesh_10_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_9_io_in_control_1_shift_pipe_b <= mesh_10_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_9_io_in_control_1_dataflow_pipe_b <= mesh_10_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_9_io_in_control_1_propagate_pipe_b <= mesh_10_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_9_io_in_control_0_shift_pipe_b <= mesh_11_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_9_io_in_control_0_dataflow_pipe_b <= mesh_11_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_9_io_in_control_0_propagate_pipe_b <= mesh_11_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_9_io_in_control_1_shift_pipe_b <= mesh_11_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_9_io_in_control_1_dataflow_pipe_b <= mesh_11_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_9_io_in_control_1_propagate_pipe_b <= mesh_11_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_9_io_in_control_0_shift_pipe_b <= mesh_12_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_9_io_in_control_0_dataflow_pipe_b <= mesh_12_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_9_io_in_control_0_propagate_pipe_b <= mesh_12_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_9_io_in_control_1_shift_pipe_b <= mesh_12_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_9_io_in_control_1_dataflow_pipe_b <= mesh_12_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_9_io_in_control_1_propagate_pipe_b <= mesh_12_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_9_io_in_control_0_shift_pipe_b <= mesh_13_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_9_io_in_control_0_dataflow_pipe_b <= mesh_13_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_9_io_in_control_0_propagate_pipe_b <= mesh_13_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_9_io_in_control_1_shift_pipe_b <= mesh_13_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_9_io_in_control_1_dataflow_pipe_b <= mesh_13_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_9_io_in_control_1_propagate_pipe_b <= mesh_13_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_9_io_in_control_0_shift_pipe_b <= mesh_14_9_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_9_io_in_control_0_dataflow_pipe_b <= mesh_14_9_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_9_io_in_control_0_propagate_pipe_b <= mesh_14_9_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_9_io_in_control_1_shift_pipe_b <= mesh_14_9_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_9_io_in_control_1_dataflow_pipe_b <= mesh_14_9_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_9_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_9_io_in_control_1_propagate_pipe_b <= mesh_14_9_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_10_io_in_control_0_shift_pipe_b <= io_in_control_10_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_10_io_in_control_0_dataflow_pipe_b <= io_in_control_10_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_10_io_in_control_0_propagate_pipe_b <= io_in_control_10_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_10_io_in_control_1_shift_pipe_b <= io_in_control_10_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_10_io_in_control_1_dataflow_pipe_b <= io_in_control_10_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_10_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_10_io_in_control_1_propagate_pipe_b <= io_in_control_10_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_10_io_in_control_0_shift_pipe_b <= mesh_0_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_10_io_in_control_0_dataflow_pipe_b <= mesh_0_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_10_io_in_control_0_propagate_pipe_b <= mesh_0_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_10_io_in_control_1_shift_pipe_b <= mesh_0_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_10_io_in_control_1_dataflow_pipe_b <= mesh_0_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_10_io_in_control_1_propagate_pipe_b <= mesh_0_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_10_io_in_control_0_shift_pipe_b <= mesh_1_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_10_io_in_control_0_dataflow_pipe_b <= mesh_1_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_10_io_in_control_0_propagate_pipe_b <= mesh_1_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_10_io_in_control_1_shift_pipe_b <= mesh_1_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_10_io_in_control_1_dataflow_pipe_b <= mesh_1_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_10_io_in_control_1_propagate_pipe_b <= mesh_1_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_10_io_in_control_0_shift_pipe_b <= mesh_2_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_10_io_in_control_0_dataflow_pipe_b <= mesh_2_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_10_io_in_control_0_propagate_pipe_b <= mesh_2_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_10_io_in_control_1_shift_pipe_b <= mesh_2_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_10_io_in_control_1_dataflow_pipe_b <= mesh_2_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_10_io_in_control_1_propagate_pipe_b <= mesh_2_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_10_io_in_control_0_shift_pipe_b <= mesh_3_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_10_io_in_control_0_dataflow_pipe_b <= mesh_3_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_10_io_in_control_0_propagate_pipe_b <= mesh_3_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_10_io_in_control_1_shift_pipe_b <= mesh_3_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_10_io_in_control_1_dataflow_pipe_b <= mesh_3_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_10_io_in_control_1_propagate_pipe_b <= mesh_3_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_10_io_in_control_0_shift_pipe_b <= mesh_4_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_10_io_in_control_0_dataflow_pipe_b <= mesh_4_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_10_io_in_control_0_propagate_pipe_b <= mesh_4_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_10_io_in_control_1_shift_pipe_b <= mesh_4_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_10_io_in_control_1_dataflow_pipe_b <= mesh_4_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_10_io_in_control_1_propagate_pipe_b <= mesh_4_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_10_io_in_control_0_shift_pipe_b <= mesh_5_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_10_io_in_control_0_dataflow_pipe_b <= mesh_5_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_10_io_in_control_0_propagate_pipe_b <= mesh_5_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_10_io_in_control_1_shift_pipe_b <= mesh_5_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_10_io_in_control_1_dataflow_pipe_b <= mesh_5_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_10_io_in_control_1_propagate_pipe_b <= mesh_5_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_10_io_in_control_0_shift_pipe_b <= mesh_6_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_10_io_in_control_0_dataflow_pipe_b <= mesh_6_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_10_io_in_control_0_propagate_pipe_b <= mesh_6_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_10_io_in_control_1_shift_pipe_b <= mesh_6_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_10_io_in_control_1_dataflow_pipe_b <= mesh_6_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_10_io_in_control_1_propagate_pipe_b <= mesh_6_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_10_io_in_control_0_shift_pipe_b <= mesh_7_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_10_io_in_control_0_dataflow_pipe_b <= mesh_7_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_10_io_in_control_0_propagate_pipe_b <= mesh_7_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_10_io_in_control_1_shift_pipe_b <= mesh_7_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_10_io_in_control_1_dataflow_pipe_b <= mesh_7_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_10_io_in_control_1_propagate_pipe_b <= mesh_7_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_10_io_in_control_0_shift_pipe_b <= mesh_8_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_10_io_in_control_0_dataflow_pipe_b <= mesh_8_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_10_io_in_control_0_propagate_pipe_b <= mesh_8_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_10_io_in_control_1_shift_pipe_b <= mesh_8_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_10_io_in_control_1_dataflow_pipe_b <= mesh_8_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_10_io_in_control_1_propagate_pipe_b <= mesh_8_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_10_io_in_control_0_shift_pipe_b <= mesh_9_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_10_io_in_control_0_dataflow_pipe_b <= mesh_9_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_10_io_in_control_0_propagate_pipe_b <= mesh_9_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_10_io_in_control_1_shift_pipe_b <= mesh_9_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_10_io_in_control_1_dataflow_pipe_b <= mesh_9_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_10_io_in_control_1_propagate_pipe_b <= mesh_9_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_10_io_in_control_0_shift_pipe_b <= mesh_10_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_10_io_in_control_0_dataflow_pipe_b <= mesh_10_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_10_io_in_control_0_propagate_pipe_b <= mesh_10_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_10_io_in_control_1_shift_pipe_b <= mesh_10_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_10_io_in_control_1_dataflow_pipe_b <= mesh_10_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_10_io_in_control_1_propagate_pipe_b <= mesh_10_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_10_io_in_control_0_shift_pipe_b <= mesh_11_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_10_io_in_control_0_dataflow_pipe_b <= mesh_11_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_10_io_in_control_0_propagate_pipe_b <= mesh_11_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_10_io_in_control_1_shift_pipe_b <= mesh_11_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_10_io_in_control_1_dataflow_pipe_b <= mesh_11_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_10_io_in_control_1_propagate_pipe_b <= mesh_11_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_10_io_in_control_0_shift_pipe_b <= mesh_12_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_10_io_in_control_0_dataflow_pipe_b <= mesh_12_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_10_io_in_control_0_propagate_pipe_b <= mesh_12_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_10_io_in_control_1_shift_pipe_b <= mesh_12_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_10_io_in_control_1_dataflow_pipe_b <= mesh_12_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_10_io_in_control_1_propagate_pipe_b <= mesh_12_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_10_io_in_control_0_shift_pipe_b <= mesh_13_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_10_io_in_control_0_dataflow_pipe_b <= mesh_13_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_10_io_in_control_0_propagate_pipe_b <= mesh_13_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_10_io_in_control_1_shift_pipe_b <= mesh_13_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_10_io_in_control_1_dataflow_pipe_b <= mesh_13_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_10_io_in_control_1_propagate_pipe_b <= mesh_13_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_10_io_in_control_0_shift_pipe_b <= mesh_14_10_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_10_io_in_control_0_dataflow_pipe_b <= mesh_14_10_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_10_io_in_control_0_propagate_pipe_b <= mesh_14_10_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_10_io_in_control_1_shift_pipe_b <= mesh_14_10_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_10_io_in_control_1_dataflow_pipe_b <= mesh_14_10_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_10_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_10_io_in_control_1_propagate_pipe_b <= mesh_14_10_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_11_io_in_control_0_shift_pipe_b <= io_in_control_11_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_11_io_in_control_0_dataflow_pipe_b <= io_in_control_11_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_11_io_in_control_0_propagate_pipe_b <= io_in_control_11_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_11_io_in_control_1_shift_pipe_b <= io_in_control_11_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_11_io_in_control_1_dataflow_pipe_b <= io_in_control_11_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_11_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_11_io_in_control_1_propagate_pipe_b <= io_in_control_11_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_11_io_in_control_0_shift_pipe_b <= mesh_0_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_11_io_in_control_0_dataflow_pipe_b <= mesh_0_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_11_io_in_control_0_propagate_pipe_b <= mesh_0_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_11_io_in_control_1_shift_pipe_b <= mesh_0_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_11_io_in_control_1_dataflow_pipe_b <= mesh_0_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_11_io_in_control_1_propagate_pipe_b <= mesh_0_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_11_io_in_control_0_shift_pipe_b <= mesh_1_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_11_io_in_control_0_dataflow_pipe_b <= mesh_1_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_11_io_in_control_0_propagate_pipe_b <= mesh_1_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_11_io_in_control_1_shift_pipe_b <= mesh_1_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_11_io_in_control_1_dataflow_pipe_b <= mesh_1_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_11_io_in_control_1_propagate_pipe_b <= mesh_1_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_11_io_in_control_0_shift_pipe_b <= mesh_2_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_11_io_in_control_0_dataflow_pipe_b <= mesh_2_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_11_io_in_control_0_propagate_pipe_b <= mesh_2_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_11_io_in_control_1_shift_pipe_b <= mesh_2_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_11_io_in_control_1_dataflow_pipe_b <= mesh_2_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_11_io_in_control_1_propagate_pipe_b <= mesh_2_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_11_io_in_control_0_shift_pipe_b <= mesh_3_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_11_io_in_control_0_dataflow_pipe_b <= mesh_3_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_11_io_in_control_0_propagate_pipe_b <= mesh_3_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_11_io_in_control_1_shift_pipe_b <= mesh_3_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_11_io_in_control_1_dataflow_pipe_b <= mesh_3_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_11_io_in_control_1_propagate_pipe_b <= mesh_3_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_11_io_in_control_0_shift_pipe_b <= mesh_4_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_11_io_in_control_0_dataflow_pipe_b <= mesh_4_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_11_io_in_control_0_propagate_pipe_b <= mesh_4_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_11_io_in_control_1_shift_pipe_b <= mesh_4_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_11_io_in_control_1_dataflow_pipe_b <= mesh_4_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_11_io_in_control_1_propagate_pipe_b <= mesh_4_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_11_io_in_control_0_shift_pipe_b <= mesh_5_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_11_io_in_control_0_dataflow_pipe_b <= mesh_5_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_11_io_in_control_0_propagate_pipe_b <= mesh_5_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_11_io_in_control_1_shift_pipe_b <= mesh_5_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_11_io_in_control_1_dataflow_pipe_b <= mesh_5_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_11_io_in_control_1_propagate_pipe_b <= mesh_5_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_11_io_in_control_0_shift_pipe_b <= mesh_6_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_11_io_in_control_0_dataflow_pipe_b <= mesh_6_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_11_io_in_control_0_propagate_pipe_b <= mesh_6_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_11_io_in_control_1_shift_pipe_b <= mesh_6_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_11_io_in_control_1_dataflow_pipe_b <= mesh_6_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_11_io_in_control_1_propagate_pipe_b <= mesh_6_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_11_io_in_control_0_shift_pipe_b <= mesh_7_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_11_io_in_control_0_dataflow_pipe_b <= mesh_7_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_11_io_in_control_0_propagate_pipe_b <= mesh_7_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_11_io_in_control_1_shift_pipe_b <= mesh_7_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_11_io_in_control_1_dataflow_pipe_b <= mesh_7_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_11_io_in_control_1_propagate_pipe_b <= mesh_7_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_11_io_in_control_0_shift_pipe_b <= mesh_8_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_11_io_in_control_0_dataflow_pipe_b <= mesh_8_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_11_io_in_control_0_propagate_pipe_b <= mesh_8_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_11_io_in_control_1_shift_pipe_b <= mesh_8_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_11_io_in_control_1_dataflow_pipe_b <= mesh_8_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_11_io_in_control_1_propagate_pipe_b <= mesh_8_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_11_io_in_control_0_shift_pipe_b <= mesh_9_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_11_io_in_control_0_dataflow_pipe_b <= mesh_9_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_11_io_in_control_0_propagate_pipe_b <= mesh_9_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_11_io_in_control_1_shift_pipe_b <= mesh_9_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_11_io_in_control_1_dataflow_pipe_b <= mesh_9_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_11_io_in_control_1_propagate_pipe_b <= mesh_9_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_11_io_in_control_0_shift_pipe_b <= mesh_10_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_11_io_in_control_0_dataflow_pipe_b <= mesh_10_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_11_io_in_control_0_propagate_pipe_b <= mesh_10_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_11_io_in_control_1_shift_pipe_b <= mesh_10_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_11_io_in_control_1_dataflow_pipe_b <= mesh_10_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_11_io_in_control_1_propagate_pipe_b <= mesh_10_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_11_io_in_control_0_shift_pipe_b <= mesh_11_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_11_io_in_control_0_dataflow_pipe_b <= mesh_11_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_11_io_in_control_0_propagate_pipe_b <= mesh_11_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_11_io_in_control_1_shift_pipe_b <= mesh_11_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_11_io_in_control_1_dataflow_pipe_b <= mesh_11_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_11_io_in_control_1_propagate_pipe_b <= mesh_11_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_11_io_in_control_0_shift_pipe_b <= mesh_12_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_11_io_in_control_0_dataflow_pipe_b <= mesh_12_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_11_io_in_control_0_propagate_pipe_b <= mesh_12_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_11_io_in_control_1_shift_pipe_b <= mesh_12_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_11_io_in_control_1_dataflow_pipe_b <= mesh_12_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_11_io_in_control_1_propagate_pipe_b <= mesh_12_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_11_io_in_control_0_shift_pipe_b <= mesh_13_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_11_io_in_control_0_dataflow_pipe_b <= mesh_13_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_11_io_in_control_0_propagate_pipe_b <= mesh_13_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_11_io_in_control_1_shift_pipe_b <= mesh_13_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_11_io_in_control_1_dataflow_pipe_b <= mesh_13_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_11_io_in_control_1_propagate_pipe_b <= mesh_13_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_11_io_in_control_0_shift_pipe_b <= mesh_14_11_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_11_io_in_control_0_dataflow_pipe_b <= mesh_14_11_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_11_io_in_control_0_propagate_pipe_b <= mesh_14_11_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_11_io_in_control_1_shift_pipe_b <= mesh_14_11_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_11_io_in_control_1_dataflow_pipe_b <= mesh_14_11_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_11_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_11_io_in_control_1_propagate_pipe_b <= mesh_14_11_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_12_io_in_control_0_shift_pipe_b <= io_in_control_12_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_12_io_in_control_0_dataflow_pipe_b <= io_in_control_12_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_12_io_in_control_0_propagate_pipe_b <= io_in_control_12_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_12_io_in_control_1_shift_pipe_b <= io_in_control_12_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_12_io_in_control_1_dataflow_pipe_b <= io_in_control_12_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_12_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_12_io_in_control_1_propagate_pipe_b <= io_in_control_12_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_12_io_in_control_0_shift_pipe_b <= mesh_0_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_12_io_in_control_0_dataflow_pipe_b <= mesh_0_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_12_io_in_control_0_propagate_pipe_b <= mesh_0_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_12_io_in_control_1_shift_pipe_b <= mesh_0_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_12_io_in_control_1_dataflow_pipe_b <= mesh_0_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_12_io_in_control_1_propagate_pipe_b <= mesh_0_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_12_io_in_control_0_shift_pipe_b <= mesh_1_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_12_io_in_control_0_dataflow_pipe_b <= mesh_1_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_12_io_in_control_0_propagate_pipe_b <= mesh_1_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_12_io_in_control_1_shift_pipe_b <= mesh_1_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_12_io_in_control_1_dataflow_pipe_b <= mesh_1_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_12_io_in_control_1_propagate_pipe_b <= mesh_1_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_12_io_in_control_0_shift_pipe_b <= mesh_2_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_12_io_in_control_0_dataflow_pipe_b <= mesh_2_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_12_io_in_control_0_propagate_pipe_b <= mesh_2_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_12_io_in_control_1_shift_pipe_b <= mesh_2_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_12_io_in_control_1_dataflow_pipe_b <= mesh_2_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_12_io_in_control_1_propagate_pipe_b <= mesh_2_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_12_io_in_control_0_shift_pipe_b <= mesh_3_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_12_io_in_control_0_dataflow_pipe_b <= mesh_3_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_12_io_in_control_0_propagate_pipe_b <= mesh_3_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_12_io_in_control_1_shift_pipe_b <= mesh_3_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_12_io_in_control_1_dataflow_pipe_b <= mesh_3_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_12_io_in_control_1_propagate_pipe_b <= mesh_3_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_12_io_in_control_0_shift_pipe_b <= mesh_4_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_12_io_in_control_0_dataflow_pipe_b <= mesh_4_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_12_io_in_control_0_propagate_pipe_b <= mesh_4_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_12_io_in_control_1_shift_pipe_b <= mesh_4_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_12_io_in_control_1_dataflow_pipe_b <= mesh_4_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_12_io_in_control_1_propagate_pipe_b <= mesh_4_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_12_io_in_control_0_shift_pipe_b <= mesh_5_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_12_io_in_control_0_dataflow_pipe_b <= mesh_5_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_12_io_in_control_0_propagate_pipe_b <= mesh_5_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_12_io_in_control_1_shift_pipe_b <= mesh_5_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_12_io_in_control_1_dataflow_pipe_b <= mesh_5_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_12_io_in_control_1_propagate_pipe_b <= mesh_5_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_12_io_in_control_0_shift_pipe_b <= mesh_6_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_12_io_in_control_0_dataflow_pipe_b <= mesh_6_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_12_io_in_control_0_propagate_pipe_b <= mesh_6_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_12_io_in_control_1_shift_pipe_b <= mesh_6_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_12_io_in_control_1_dataflow_pipe_b <= mesh_6_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_12_io_in_control_1_propagate_pipe_b <= mesh_6_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_12_io_in_control_0_shift_pipe_b <= mesh_7_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_12_io_in_control_0_dataflow_pipe_b <= mesh_7_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_12_io_in_control_0_propagate_pipe_b <= mesh_7_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_12_io_in_control_1_shift_pipe_b <= mesh_7_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_12_io_in_control_1_dataflow_pipe_b <= mesh_7_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_12_io_in_control_1_propagate_pipe_b <= mesh_7_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_12_io_in_control_0_shift_pipe_b <= mesh_8_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_12_io_in_control_0_dataflow_pipe_b <= mesh_8_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_12_io_in_control_0_propagate_pipe_b <= mesh_8_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_12_io_in_control_1_shift_pipe_b <= mesh_8_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_12_io_in_control_1_dataflow_pipe_b <= mesh_8_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_12_io_in_control_1_propagate_pipe_b <= mesh_8_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_12_io_in_control_0_shift_pipe_b <= mesh_9_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_12_io_in_control_0_dataflow_pipe_b <= mesh_9_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_12_io_in_control_0_propagate_pipe_b <= mesh_9_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_12_io_in_control_1_shift_pipe_b <= mesh_9_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_12_io_in_control_1_dataflow_pipe_b <= mesh_9_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_12_io_in_control_1_propagate_pipe_b <= mesh_9_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_12_io_in_control_0_shift_pipe_b <= mesh_10_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_12_io_in_control_0_dataflow_pipe_b <= mesh_10_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_12_io_in_control_0_propagate_pipe_b <= mesh_10_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_12_io_in_control_1_shift_pipe_b <= mesh_10_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_12_io_in_control_1_dataflow_pipe_b <= mesh_10_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_12_io_in_control_1_propagate_pipe_b <= mesh_10_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_12_io_in_control_0_shift_pipe_b <= mesh_11_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_12_io_in_control_0_dataflow_pipe_b <= mesh_11_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_12_io_in_control_0_propagate_pipe_b <= mesh_11_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_12_io_in_control_1_shift_pipe_b <= mesh_11_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_12_io_in_control_1_dataflow_pipe_b <= mesh_11_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_12_io_in_control_1_propagate_pipe_b <= mesh_11_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_12_io_in_control_0_shift_pipe_b <= mesh_12_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_12_io_in_control_0_dataflow_pipe_b <= mesh_12_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_12_io_in_control_0_propagate_pipe_b <= mesh_12_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_12_io_in_control_1_shift_pipe_b <= mesh_12_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_12_io_in_control_1_dataflow_pipe_b <= mesh_12_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_12_io_in_control_1_propagate_pipe_b <= mesh_12_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_12_io_in_control_0_shift_pipe_b <= mesh_13_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_12_io_in_control_0_dataflow_pipe_b <= mesh_13_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_12_io_in_control_0_propagate_pipe_b <= mesh_13_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_12_io_in_control_1_shift_pipe_b <= mesh_13_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_12_io_in_control_1_dataflow_pipe_b <= mesh_13_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_12_io_in_control_1_propagate_pipe_b <= mesh_13_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_12_io_in_control_0_shift_pipe_b <= mesh_14_12_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_12_io_in_control_0_dataflow_pipe_b <= mesh_14_12_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_12_io_in_control_0_propagate_pipe_b <= mesh_14_12_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_12_io_in_control_1_shift_pipe_b <= mesh_14_12_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_12_io_in_control_1_dataflow_pipe_b <= mesh_14_12_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_12_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_12_io_in_control_1_propagate_pipe_b <= mesh_14_12_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_13_io_in_control_0_shift_pipe_b <= io_in_control_13_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_13_io_in_control_0_dataflow_pipe_b <= io_in_control_13_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_13_io_in_control_0_propagate_pipe_b <= io_in_control_13_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_13_io_in_control_1_shift_pipe_b <= io_in_control_13_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_13_io_in_control_1_dataflow_pipe_b <= io_in_control_13_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_13_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_13_io_in_control_1_propagate_pipe_b <= io_in_control_13_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_13_io_in_control_0_shift_pipe_b <= mesh_0_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_13_io_in_control_0_dataflow_pipe_b <= mesh_0_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_13_io_in_control_0_propagate_pipe_b <= mesh_0_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_13_io_in_control_1_shift_pipe_b <= mesh_0_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_13_io_in_control_1_dataflow_pipe_b <= mesh_0_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_13_io_in_control_1_propagate_pipe_b <= mesh_0_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_13_io_in_control_0_shift_pipe_b <= mesh_1_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_13_io_in_control_0_dataflow_pipe_b <= mesh_1_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_13_io_in_control_0_propagate_pipe_b <= mesh_1_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_13_io_in_control_1_shift_pipe_b <= mesh_1_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_13_io_in_control_1_dataflow_pipe_b <= mesh_1_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_13_io_in_control_1_propagate_pipe_b <= mesh_1_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_13_io_in_control_0_shift_pipe_b <= mesh_2_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_13_io_in_control_0_dataflow_pipe_b <= mesh_2_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_13_io_in_control_0_propagate_pipe_b <= mesh_2_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_13_io_in_control_1_shift_pipe_b <= mesh_2_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_13_io_in_control_1_dataflow_pipe_b <= mesh_2_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_13_io_in_control_1_propagate_pipe_b <= mesh_2_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_13_io_in_control_0_shift_pipe_b <= mesh_3_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_13_io_in_control_0_dataflow_pipe_b <= mesh_3_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_13_io_in_control_0_propagate_pipe_b <= mesh_3_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_13_io_in_control_1_shift_pipe_b <= mesh_3_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_13_io_in_control_1_dataflow_pipe_b <= mesh_3_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_13_io_in_control_1_propagate_pipe_b <= mesh_3_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_13_io_in_control_0_shift_pipe_b <= mesh_4_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_13_io_in_control_0_dataflow_pipe_b <= mesh_4_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_13_io_in_control_0_propagate_pipe_b <= mesh_4_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_13_io_in_control_1_shift_pipe_b <= mesh_4_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_13_io_in_control_1_dataflow_pipe_b <= mesh_4_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_13_io_in_control_1_propagate_pipe_b <= mesh_4_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_13_io_in_control_0_shift_pipe_b <= mesh_5_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_13_io_in_control_0_dataflow_pipe_b <= mesh_5_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_13_io_in_control_0_propagate_pipe_b <= mesh_5_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_13_io_in_control_1_shift_pipe_b <= mesh_5_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_13_io_in_control_1_dataflow_pipe_b <= mesh_5_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_13_io_in_control_1_propagate_pipe_b <= mesh_5_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_13_io_in_control_0_shift_pipe_b <= mesh_6_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_13_io_in_control_0_dataflow_pipe_b <= mesh_6_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_13_io_in_control_0_propagate_pipe_b <= mesh_6_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_13_io_in_control_1_shift_pipe_b <= mesh_6_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_13_io_in_control_1_dataflow_pipe_b <= mesh_6_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_13_io_in_control_1_propagate_pipe_b <= mesh_6_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_13_io_in_control_0_shift_pipe_b <= mesh_7_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_13_io_in_control_0_dataflow_pipe_b <= mesh_7_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_13_io_in_control_0_propagate_pipe_b <= mesh_7_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_13_io_in_control_1_shift_pipe_b <= mesh_7_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_13_io_in_control_1_dataflow_pipe_b <= mesh_7_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_13_io_in_control_1_propagate_pipe_b <= mesh_7_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_13_io_in_control_0_shift_pipe_b <= mesh_8_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_13_io_in_control_0_dataflow_pipe_b <= mesh_8_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_13_io_in_control_0_propagate_pipe_b <= mesh_8_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_13_io_in_control_1_shift_pipe_b <= mesh_8_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_13_io_in_control_1_dataflow_pipe_b <= mesh_8_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_13_io_in_control_1_propagate_pipe_b <= mesh_8_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_13_io_in_control_0_shift_pipe_b <= mesh_9_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_13_io_in_control_0_dataflow_pipe_b <= mesh_9_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_13_io_in_control_0_propagate_pipe_b <= mesh_9_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_13_io_in_control_1_shift_pipe_b <= mesh_9_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_13_io_in_control_1_dataflow_pipe_b <= mesh_9_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_13_io_in_control_1_propagate_pipe_b <= mesh_9_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_13_io_in_control_0_shift_pipe_b <= mesh_10_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_13_io_in_control_0_dataflow_pipe_b <= mesh_10_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_13_io_in_control_0_propagate_pipe_b <= mesh_10_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_13_io_in_control_1_shift_pipe_b <= mesh_10_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_13_io_in_control_1_dataflow_pipe_b <= mesh_10_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_13_io_in_control_1_propagate_pipe_b <= mesh_10_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_13_io_in_control_0_shift_pipe_b <= mesh_11_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_13_io_in_control_0_dataflow_pipe_b <= mesh_11_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_13_io_in_control_0_propagate_pipe_b <= mesh_11_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_13_io_in_control_1_shift_pipe_b <= mesh_11_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_13_io_in_control_1_dataflow_pipe_b <= mesh_11_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_13_io_in_control_1_propagate_pipe_b <= mesh_11_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_13_io_in_control_0_shift_pipe_b <= mesh_12_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_13_io_in_control_0_dataflow_pipe_b <= mesh_12_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_13_io_in_control_0_propagate_pipe_b <= mesh_12_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_13_io_in_control_1_shift_pipe_b <= mesh_12_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_13_io_in_control_1_dataflow_pipe_b <= mesh_12_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_13_io_in_control_1_propagate_pipe_b <= mesh_12_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_13_io_in_control_0_shift_pipe_b <= mesh_13_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_13_io_in_control_0_dataflow_pipe_b <= mesh_13_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_13_io_in_control_0_propagate_pipe_b <= mesh_13_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_13_io_in_control_1_shift_pipe_b <= mesh_13_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_13_io_in_control_1_dataflow_pipe_b <= mesh_13_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_13_io_in_control_1_propagate_pipe_b <= mesh_13_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_13_io_in_control_0_shift_pipe_b <= mesh_14_13_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_13_io_in_control_0_dataflow_pipe_b <= mesh_14_13_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_13_io_in_control_0_propagate_pipe_b <= mesh_14_13_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_13_io_in_control_1_shift_pipe_b <= mesh_14_13_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_13_io_in_control_1_dataflow_pipe_b <= mesh_14_13_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_13_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_13_io_in_control_1_propagate_pipe_b <= mesh_14_13_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_14_io_in_control_0_shift_pipe_b <= io_in_control_14_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_14_io_in_control_0_dataflow_pipe_b <= io_in_control_14_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_14_io_in_control_0_propagate_pipe_b <= io_in_control_14_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_14_io_in_control_1_shift_pipe_b <= io_in_control_14_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_14_io_in_control_1_dataflow_pipe_b <= io_in_control_14_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_14_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_14_io_in_control_1_propagate_pipe_b <= io_in_control_14_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_14_io_in_control_0_shift_pipe_b <= mesh_0_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_14_io_in_control_0_dataflow_pipe_b <= mesh_0_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_14_io_in_control_0_propagate_pipe_b <= mesh_0_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_14_io_in_control_1_shift_pipe_b <= mesh_0_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_14_io_in_control_1_dataflow_pipe_b <= mesh_0_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_14_io_in_control_1_propagate_pipe_b <= mesh_0_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_14_io_in_control_0_shift_pipe_b <= mesh_1_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_14_io_in_control_0_dataflow_pipe_b <= mesh_1_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_14_io_in_control_0_propagate_pipe_b <= mesh_1_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_14_io_in_control_1_shift_pipe_b <= mesh_1_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_14_io_in_control_1_dataflow_pipe_b <= mesh_1_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_14_io_in_control_1_propagate_pipe_b <= mesh_1_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_14_io_in_control_0_shift_pipe_b <= mesh_2_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_14_io_in_control_0_dataflow_pipe_b <= mesh_2_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_14_io_in_control_0_propagate_pipe_b <= mesh_2_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_14_io_in_control_1_shift_pipe_b <= mesh_2_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_14_io_in_control_1_dataflow_pipe_b <= mesh_2_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_14_io_in_control_1_propagate_pipe_b <= mesh_2_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_14_io_in_control_0_shift_pipe_b <= mesh_3_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_14_io_in_control_0_dataflow_pipe_b <= mesh_3_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_14_io_in_control_0_propagate_pipe_b <= mesh_3_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_14_io_in_control_1_shift_pipe_b <= mesh_3_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_14_io_in_control_1_dataflow_pipe_b <= mesh_3_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_14_io_in_control_1_propagate_pipe_b <= mesh_3_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_14_io_in_control_0_shift_pipe_b <= mesh_4_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_14_io_in_control_0_dataflow_pipe_b <= mesh_4_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_14_io_in_control_0_propagate_pipe_b <= mesh_4_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_14_io_in_control_1_shift_pipe_b <= mesh_4_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_14_io_in_control_1_dataflow_pipe_b <= mesh_4_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_14_io_in_control_1_propagate_pipe_b <= mesh_4_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_14_io_in_control_0_shift_pipe_b <= mesh_5_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_14_io_in_control_0_dataflow_pipe_b <= mesh_5_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_14_io_in_control_0_propagate_pipe_b <= mesh_5_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_14_io_in_control_1_shift_pipe_b <= mesh_5_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_14_io_in_control_1_dataflow_pipe_b <= mesh_5_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_14_io_in_control_1_propagate_pipe_b <= mesh_5_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_14_io_in_control_0_shift_pipe_b <= mesh_6_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_14_io_in_control_0_dataflow_pipe_b <= mesh_6_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_14_io_in_control_0_propagate_pipe_b <= mesh_6_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_14_io_in_control_1_shift_pipe_b <= mesh_6_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_14_io_in_control_1_dataflow_pipe_b <= mesh_6_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_14_io_in_control_1_propagate_pipe_b <= mesh_6_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_14_io_in_control_0_shift_pipe_b <= mesh_7_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_14_io_in_control_0_dataflow_pipe_b <= mesh_7_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_14_io_in_control_0_propagate_pipe_b <= mesh_7_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_14_io_in_control_1_shift_pipe_b <= mesh_7_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_14_io_in_control_1_dataflow_pipe_b <= mesh_7_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_14_io_in_control_1_propagate_pipe_b <= mesh_7_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_14_io_in_control_0_shift_pipe_b <= mesh_8_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_14_io_in_control_0_dataflow_pipe_b <= mesh_8_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_14_io_in_control_0_propagate_pipe_b <= mesh_8_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_14_io_in_control_1_shift_pipe_b <= mesh_8_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_14_io_in_control_1_dataflow_pipe_b <= mesh_8_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_14_io_in_control_1_propagate_pipe_b <= mesh_8_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_14_io_in_control_0_shift_pipe_b <= mesh_9_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_14_io_in_control_0_dataflow_pipe_b <= mesh_9_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_14_io_in_control_0_propagate_pipe_b <= mesh_9_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_14_io_in_control_1_shift_pipe_b <= mesh_9_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_14_io_in_control_1_dataflow_pipe_b <= mesh_9_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_14_io_in_control_1_propagate_pipe_b <= mesh_9_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_14_io_in_control_0_shift_pipe_b <= mesh_10_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_14_io_in_control_0_dataflow_pipe_b <= mesh_10_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_14_io_in_control_0_propagate_pipe_b <= mesh_10_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_14_io_in_control_1_shift_pipe_b <= mesh_10_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_14_io_in_control_1_dataflow_pipe_b <= mesh_10_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_14_io_in_control_1_propagate_pipe_b <= mesh_10_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_14_io_in_control_0_shift_pipe_b <= mesh_11_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_14_io_in_control_0_dataflow_pipe_b <= mesh_11_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_14_io_in_control_0_propagate_pipe_b <= mesh_11_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_14_io_in_control_1_shift_pipe_b <= mesh_11_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_14_io_in_control_1_dataflow_pipe_b <= mesh_11_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_14_io_in_control_1_propagate_pipe_b <= mesh_11_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_14_io_in_control_0_shift_pipe_b <= mesh_12_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_14_io_in_control_0_dataflow_pipe_b <= mesh_12_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_14_io_in_control_0_propagate_pipe_b <= mesh_12_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_14_io_in_control_1_shift_pipe_b <= mesh_12_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_14_io_in_control_1_dataflow_pipe_b <= mesh_12_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_14_io_in_control_1_propagate_pipe_b <= mesh_12_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_14_io_in_control_0_shift_pipe_b <= mesh_13_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_14_io_in_control_0_dataflow_pipe_b <= mesh_13_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_14_io_in_control_0_propagate_pipe_b <= mesh_13_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_14_io_in_control_1_shift_pipe_b <= mesh_13_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_14_io_in_control_1_dataflow_pipe_b <= mesh_13_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_14_io_in_control_1_propagate_pipe_b <= mesh_13_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_14_io_in_control_0_shift_pipe_b <= mesh_14_14_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_14_io_in_control_0_dataflow_pipe_b <= mesh_14_14_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_14_io_in_control_0_propagate_pipe_b <= mesh_14_14_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_14_io_in_control_1_shift_pipe_b <= mesh_14_14_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_14_io_in_control_1_dataflow_pipe_b <= mesh_14_14_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_14_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_14_io_in_control_1_propagate_pipe_b <= mesh_14_14_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_15_io_in_control_0_shift_pipe_b <= io_in_control_15_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_15_io_in_control_0_dataflow_pipe_b <= io_in_control_15_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_15_io_in_control_0_propagate_pipe_b <= io_in_control_15_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_15_io_in_control_1_shift_pipe_b <= io_in_control_15_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_15_io_in_control_1_dataflow_pipe_b <= io_in_control_15_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (io_in_valid_15_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_0_15_io_in_control_1_propagate_pipe_b <= io_in_control_15_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_15_io_in_control_0_shift_pipe_b <= mesh_0_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_15_io_in_control_0_dataflow_pipe_b <= mesh_0_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_15_io_in_control_0_propagate_pipe_b <= mesh_0_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_15_io_in_control_1_shift_pipe_b <= mesh_0_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_15_io_in_control_1_dataflow_pipe_b <= mesh_0_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_0_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_1_15_io_in_control_1_propagate_pipe_b <= mesh_0_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_15_io_in_control_0_shift_pipe_b <= mesh_1_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_15_io_in_control_0_dataflow_pipe_b <= mesh_1_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_15_io_in_control_0_propagate_pipe_b <= mesh_1_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_15_io_in_control_1_shift_pipe_b <= mesh_1_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_15_io_in_control_1_dataflow_pipe_b <= mesh_1_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_1_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_2_15_io_in_control_1_propagate_pipe_b <= mesh_1_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_15_io_in_control_0_shift_pipe_b <= mesh_2_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_15_io_in_control_0_dataflow_pipe_b <= mesh_2_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_15_io_in_control_0_propagate_pipe_b <= mesh_2_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_15_io_in_control_1_shift_pipe_b <= mesh_2_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_15_io_in_control_1_dataflow_pipe_b <= mesh_2_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_2_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_3_15_io_in_control_1_propagate_pipe_b <= mesh_2_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_15_io_in_control_0_shift_pipe_b <= mesh_3_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_15_io_in_control_0_dataflow_pipe_b <= mesh_3_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_15_io_in_control_0_propagate_pipe_b <= mesh_3_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_15_io_in_control_1_shift_pipe_b <= mesh_3_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_15_io_in_control_1_dataflow_pipe_b <= mesh_3_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_3_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_4_15_io_in_control_1_propagate_pipe_b <= mesh_3_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_15_io_in_control_0_shift_pipe_b <= mesh_4_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_15_io_in_control_0_dataflow_pipe_b <= mesh_4_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_15_io_in_control_0_propagate_pipe_b <= mesh_4_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_15_io_in_control_1_shift_pipe_b <= mesh_4_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_15_io_in_control_1_dataflow_pipe_b <= mesh_4_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_4_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_5_15_io_in_control_1_propagate_pipe_b <= mesh_4_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_15_io_in_control_0_shift_pipe_b <= mesh_5_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_15_io_in_control_0_dataflow_pipe_b <= mesh_5_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_15_io_in_control_0_propagate_pipe_b <= mesh_5_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_15_io_in_control_1_shift_pipe_b <= mesh_5_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_15_io_in_control_1_dataflow_pipe_b <= mesh_5_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_5_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_6_15_io_in_control_1_propagate_pipe_b <= mesh_5_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_15_io_in_control_0_shift_pipe_b <= mesh_6_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_15_io_in_control_0_dataflow_pipe_b <= mesh_6_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_15_io_in_control_0_propagate_pipe_b <= mesh_6_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_15_io_in_control_1_shift_pipe_b <= mesh_6_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_15_io_in_control_1_dataflow_pipe_b <= mesh_6_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_6_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_7_15_io_in_control_1_propagate_pipe_b <= mesh_6_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_15_io_in_control_0_shift_pipe_b <= mesh_7_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_15_io_in_control_0_dataflow_pipe_b <= mesh_7_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_15_io_in_control_0_propagate_pipe_b <= mesh_7_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_15_io_in_control_1_shift_pipe_b <= mesh_7_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_15_io_in_control_1_dataflow_pipe_b <= mesh_7_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_7_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_8_15_io_in_control_1_propagate_pipe_b <= mesh_7_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_15_io_in_control_0_shift_pipe_b <= mesh_8_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_15_io_in_control_0_dataflow_pipe_b <= mesh_8_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_15_io_in_control_0_propagate_pipe_b <= mesh_8_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_15_io_in_control_1_shift_pipe_b <= mesh_8_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_15_io_in_control_1_dataflow_pipe_b <= mesh_8_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_8_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_9_15_io_in_control_1_propagate_pipe_b <= mesh_8_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_15_io_in_control_0_shift_pipe_b <= mesh_9_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_15_io_in_control_0_dataflow_pipe_b <= mesh_9_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_15_io_in_control_0_propagate_pipe_b <= mesh_9_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_15_io_in_control_1_shift_pipe_b <= mesh_9_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_15_io_in_control_1_dataflow_pipe_b <= mesh_9_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_9_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_10_15_io_in_control_1_propagate_pipe_b <= mesh_9_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_15_io_in_control_0_shift_pipe_b <= mesh_10_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_15_io_in_control_0_dataflow_pipe_b <= mesh_10_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_15_io_in_control_0_propagate_pipe_b <= mesh_10_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_15_io_in_control_1_shift_pipe_b <= mesh_10_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_15_io_in_control_1_dataflow_pipe_b <= mesh_10_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_10_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_11_15_io_in_control_1_propagate_pipe_b <= mesh_10_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_15_io_in_control_0_shift_pipe_b <= mesh_11_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_15_io_in_control_0_dataflow_pipe_b <= mesh_11_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_15_io_in_control_0_propagate_pipe_b <= mesh_11_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_15_io_in_control_1_shift_pipe_b <= mesh_11_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_15_io_in_control_1_dataflow_pipe_b <= mesh_11_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_11_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_12_15_io_in_control_1_propagate_pipe_b <= mesh_11_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_15_io_in_control_0_shift_pipe_b <= mesh_12_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_15_io_in_control_0_dataflow_pipe_b <= mesh_12_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_15_io_in_control_0_propagate_pipe_b <= mesh_12_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_15_io_in_control_1_shift_pipe_b <= mesh_12_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_15_io_in_control_1_dataflow_pipe_b <= mesh_12_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_12_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_13_15_io_in_control_1_propagate_pipe_b <= mesh_12_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_15_io_in_control_0_shift_pipe_b <= mesh_13_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_15_io_in_control_0_dataflow_pipe_b <= mesh_13_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_15_io_in_control_0_propagate_pipe_b <= mesh_13_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_15_io_in_control_1_shift_pipe_b <= mesh_13_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_15_io_in_control_1_dataflow_pipe_b <= mesh_13_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_13_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_14_15_io_in_control_1_propagate_pipe_b <= mesh_13_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_15_io_in_control_0_shift_pipe_b <= mesh_14_15_io_out_control_0_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_15_io_in_control_0_dataflow_pipe_b <= mesh_14_15_io_out_control_0_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_0) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_15_io_in_control_0_propagate_pipe_b <= mesh_14_15_io_out_control_0_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_15_io_in_control_1_shift_pipe_b <= mesh_14_15_io_out_control_1_shift; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_15_io_in_control_1_dataflow_pipe_b <= mesh_14_15_io_out_control_1_dataflow; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    if (mesh_14_15_io_out_valid_1) begin // @[src/main/scala/chisel3/util/Valid.scala 135:26]
      mesh_15_15_io_in_control_1_propagate_pipe_b <= mesh_14_15_io_out_control_1_propagate; // @[src/main/scala/chisel3/util/Valid.scala 135:26]
    end
    r_256_0 <= io_in_valid_0_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_256_1 <= io_in_valid_0_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_257_0 <= mesh_0_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_257_1 <= mesh_0_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_258_0 <= mesh_1_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_258_1 <= mesh_1_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_259_0 <= mesh_2_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_259_1 <= mesh_2_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_260_0 <= mesh_3_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_260_1 <= mesh_3_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_261_0 <= mesh_4_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_261_1 <= mesh_4_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_262_0 <= mesh_5_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_262_1 <= mesh_5_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_263_0 <= mesh_6_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_263_1 <= mesh_6_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_264_0 <= mesh_7_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_264_1 <= mesh_7_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_265_0 <= mesh_8_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_265_1 <= mesh_8_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_266_0 <= mesh_9_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_266_1 <= mesh_9_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_267_0 <= mesh_10_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_267_1 <= mesh_10_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_268_0 <= mesh_11_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_268_1 <= mesh_11_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_269_0 <= mesh_12_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_269_1 <= mesh_12_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_270_0 <= mesh_13_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_270_1 <= mesh_13_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_271_0 <= mesh_14_0_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_271_1 <= mesh_14_0_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_272_0 <= io_in_valid_1_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_272_1 <= io_in_valid_1_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_273_0 <= mesh_0_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_273_1 <= mesh_0_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_274_0 <= mesh_1_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_274_1 <= mesh_1_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_275_0 <= mesh_2_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_275_1 <= mesh_2_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_276_0 <= mesh_3_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_276_1 <= mesh_3_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_277_0 <= mesh_4_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_277_1 <= mesh_4_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_278_0 <= mesh_5_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_278_1 <= mesh_5_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_279_0 <= mesh_6_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_279_1 <= mesh_6_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_280_0 <= mesh_7_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_280_1 <= mesh_7_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_281_0 <= mesh_8_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_281_1 <= mesh_8_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_282_0 <= mesh_9_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_282_1 <= mesh_9_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_283_0 <= mesh_10_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_283_1 <= mesh_10_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_284_0 <= mesh_11_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_284_1 <= mesh_11_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_285_0 <= mesh_12_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_285_1 <= mesh_12_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_286_0 <= mesh_13_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_286_1 <= mesh_13_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_287_0 <= mesh_14_1_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_287_1 <= mesh_14_1_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_288_0 <= io_in_valid_2_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_288_1 <= io_in_valid_2_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_289_0 <= mesh_0_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_289_1 <= mesh_0_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_290_0 <= mesh_1_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_290_1 <= mesh_1_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_291_0 <= mesh_2_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_291_1 <= mesh_2_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_292_0 <= mesh_3_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_292_1 <= mesh_3_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_293_0 <= mesh_4_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_293_1 <= mesh_4_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_294_0 <= mesh_5_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_294_1 <= mesh_5_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_295_0 <= mesh_6_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_295_1 <= mesh_6_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_296_0 <= mesh_7_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_296_1 <= mesh_7_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_297_0 <= mesh_8_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_297_1 <= mesh_8_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_298_0 <= mesh_9_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_298_1 <= mesh_9_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_299_0 <= mesh_10_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_299_1 <= mesh_10_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_300_0 <= mesh_11_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_300_1 <= mesh_11_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_301_0 <= mesh_12_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_301_1 <= mesh_12_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_302_0 <= mesh_13_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_302_1 <= mesh_13_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_303_0 <= mesh_14_2_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_303_1 <= mesh_14_2_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_304_0 <= io_in_valid_3_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_304_1 <= io_in_valid_3_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_305_0 <= mesh_0_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_305_1 <= mesh_0_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_306_0 <= mesh_1_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_306_1 <= mesh_1_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_307_0 <= mesh_2_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_307_1 <= mesh_2_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_308_0 <= mesh_3_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_308_1 <= mesh_3_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_309_0 <= mesh_4_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_309_1 <= mesh_4_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_310_0 <= mesh_5_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_310_1 <= mesh_5_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_311_0 <= mesh_6_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_311_1 <= mesh_6_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_312_0 <= mesh_7_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_312_1 <= mesh_7_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_313_0 <= mesh_8_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_313_1 <= mesh_8_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_314_0 <= mesh_9_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_314_1 <= mesh_9_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_315_0 <= mesh_10_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_315_1 <= mesh_10_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_316_0 <= mesh_11_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_316_1 <= mesh_11_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_317_0 <= mesh_12_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_317_1 <= mesh_12_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_318_0 <= mesh_13_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_318_1 <= mesh_13_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_319_0 <= mesh_14_3_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_319_1 <= mesh_14_3_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_320_0 <= io_in_valid_4_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_320_1 <= io_in_valid_4_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_321_0 <= mesh_0_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_321_1 <= mesh_0_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_322_0 <= mesh_1_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_322_1 <= mesh_1_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_323_0 <= mesh_2_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_323_1 <= mesh_2_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_324_0 <= mesh_3_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_324_1 <= mesh_3_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_325_0 <= mesh_4_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_325_1 <= mesh_4_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_326_0 <= mesh_5_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_326_1 <= mesh_5_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_327_0 <= mesh_6_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_327_1 <= mesh_6_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_328_0 <= mesh_7_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_328_1 <= mesh_7_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_329_0 <= mesh_8_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_329_1 <= mesh_8_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_330_0 <= mesh_9_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_330_1 <= mesh_9_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_331_0 <= mesh_10_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_331_1 <= mesh_10_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_332_0 <= mesh_11_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_332_1 <= mesh_11_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_333_0 <= mesh_12_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_333_1 <= mesh_12_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_334_0 <= mesh_13_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_334_1 <= mesh_13_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_335_0 <= mesh_14_4_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_335_1 <= mesh_14_4_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_336_0 <= io_in_valid_5_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_336_1 <= io_in_valid_5_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_337_0 <= mesh_0_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_337_1 <= mesh_0_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_338_0 <= mesh_1_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_338_1 <= mesh_1_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_339_0 <= mesh_2_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_339_1 <= mesh_2_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_340_0 <= mesh_3_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_340_1 <= mesh_3_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_341_0 <= mesh_4_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_341_1 <= mesh_4_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_342_0 <= mesh_5_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_342_1 <= mesh_5_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_343_0 <= mesh_6_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_343_1 <= mesh_6_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_344_0 <= mesh_7_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_344_1 <= mesh_7_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_345_0 <= mesh_8_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_345_1 <= mesh_8_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_346_0 <= mesh_9_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_346_1 <= mesh_9_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_347_0 <= mesh_10_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_347_1 <= mesh_10_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_348_0 <= mesh_11_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_348_1 <= mesh_11_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_349_0 <= mesh_12_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_349_1 <= mesh_12_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_350_0 <= mesh_13_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_350_1 <= mesh_13_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_351_0 <= mesh_14_5_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_351_1 <= mesh_14_5_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_352_0 <= io_in_valid_6_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_352_1 <= io_in_valid_6_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_353_0 <= mesh_0_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_353_1 <= mesh_0_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_354_0 <= mesh_1_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_354_1 <= mesh_1_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_355_0 <= mesh_2_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_355_1 <= mesh_2_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_356_0 <= mesh_3_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_356_1 <= mesh_3_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_357_0 <= mesh_4_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_357_1 <= mesh_4_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_358_0 <= mesh_5_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_358_1 <= mesh_5_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_359_0 <= mesh_6_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_359_1 <= mesh_6_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_360_0 <= mesh_7_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_360_1 <= mesh_7_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_361_0 <= mesh_8_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_361_1 <= mesh_8_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_362_0 <= mesh_9_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_362_1 <= mesh_9_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_363_0 <= mesh_10_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_363_1 <= mesh_10_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_364_0 <= mesh_11_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_364_1 <= mesh_11_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_365_0 <= mesh_12_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_365_1 <= mesh_12_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_366_0 <= mesh_13_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_366_1 <= mesh_13_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_367_0 <= mesh_14_6_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_367_1 <= mesh_14_6_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_368_0 <= io_in_valid_7_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_368_1 <= io_in_valid_7_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_369_0 <= mesh_0_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_369_1 <= mesh_0_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_370_0 <= mesh_1_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_370_1 <= mesh_1_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_371_0 <= mesh_2_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_371_1 <= mesh_2_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_372_0 <= mesh_3_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_372_1 <= mesh_3_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_373_0 <= mesh_4_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_373_1 <= mesh_4_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_374_0 <= mesh_5_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_374_1 <= mesh_5_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_375_0 <= mesh_6_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_375_1 <= mesh_6_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_376_0 <= mesh_7_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_376_1 <= mesh_7_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_377_0 <= mesh_8_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_377_1 <= mesh_8_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_378_0 <= mesh_9_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_378_1 <= mesh_9_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_379_0 <= mesh_10_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_379_1 <= mesh_10_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_380_0 <= mesh_11_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_380_1 <= mesh_11_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_381_0 <= mesh_12_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_381_1 <= mesh_12_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_382_0 <= mesh_13_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_382_1 <= mesh_13_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_383_0 <= mesh_14_7_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_383_1 <= mesh_14_7_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_384_0 <= io_in_valid_8_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_384_1 <= io_in_valid_8_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_385_0 <= mesh_0_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_385_1 <= mesh_0_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_386_0 <= mesh_1_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_386_1 <= mesh_1_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_387_0 <= mesh_2_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_387_1 <= mesh_2_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_388_0 <= mesh_3_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_388_1 <= mesh_3_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_389_0 <= mesh_4_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_389_1 <= mesh_4_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_390_0 <= mesh_5_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_390_1 <= mesh_5_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_391_0 <= mesh_6_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_391_1 <= mesh_6_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_392_0 <= mesh_7_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_392_1 <= mesh_7_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_393_0 <= mesh_8_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_393_1 <= mesh_8_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_394_0 <= mesh_9_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_394_1 <= mesh_9_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_395_0 <= mesh_10_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_395_1 <= mesh_10_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_396_0 <= mesh_11_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_396_1 <= mesh_11_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_397_0 <= mesh_12_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_397_1 <= mesh_12_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_398_0 <= mesh_13_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_398_1 <= mesh_13_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_399_0 <= mesh_14_8_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_399_1 <= mesh_14_8_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_400_0 <= io_in_valid_9_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_400_1 <= io_in_valid_9_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_401_0 <= mesh_0_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_401_1 <= mesh_0_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_402_0 <= mesh_1_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_402_1 <= mesh_1_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_403_0 <= mesh_2_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_403_1 <= mesh_2_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_404_0 <= mesh_3_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_404_1 <= mesh_3_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_405_0 <= mesh_4_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_405_1 <= mesh_4_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_406_0 <= mesh_5_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_406_1 <= mesh_5_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_407_0 <= mesh_6_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_407_1 <= mesh_6_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_408_0 <= mesh_7_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_408_1 <= mesh_7_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_409_0 <= mesh_8_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_409_1 <= mesh_8_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_410_0 <= mesh_9_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_410_1 <= mesh_9_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_411_0 <= mesh_10_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_411_1 <= mesh_10_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_412_0 <= mesh_11_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_412_1 <= mesh_11_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_413_0 <= mesh_12_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_413_1 <= mesh_12_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_414_0 <= mesh_13_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_414_1 <= mesh_13_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_415_0 <= mesh_14_9_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_415_1 <= mesh_14_9_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_416_0 <= io_in_valid_10_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_416_1 <= io_in_valid_10_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_417_0 <= mesh_0_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_417_1 <= mesh_0_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_418_0 <= mesh_1_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_418_1 <= mesh_1_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_419_0 <= mesh_2_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_419_1 <= mesh_2_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_420_0 <= mesh_3_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_420_1 <= mesh_3_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_421_0 <= mesh_4_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_421_1 <= mesh_4_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_422_0 <= mesh_5_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_422_1 <= mesh_5_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_423_0 <= mesh_6_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_423_1 <= mesh_6_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_424_0 <= mesh_7_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_424_1 <= mesh_7_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_425_0 <= mesh_8_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_425_1 <= mesh_8_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_426_0 <= mesh_9_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_426_1 <= mesh_9_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_427_0 <= mesh_10_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_427_1 <= mesh_10_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_428_0 <= mesh_11_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_428_1 <= mesh_11_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_429_0 <= mesh_12_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_429_1 <= mesh_12_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_430_0 <= mesh_13_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_430_1 <= mesh_13_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_431_0 <= mesh_14_10_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_431_1 <= mesh_14_10_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_432_0 <= io_in_valid_11_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_432_1 <= io_in_valid_11_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_433_0 <= mesh_0_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_433_1 <= mesh_0_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_434_0 <= mesh_1_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_434_1 <= mesh_1_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_435_0 <= mesh_2_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_435_1 <= mesh_2_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_436_0 <= mesh_3_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_436_1 <= mesh_3_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_437_0 <= mesh_4_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_437_1 <= mesh_4_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_438_0 <= mesh_5_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_438_1 <= mesh_5_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_439_0 <= mesh_6_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_439_1 <= mesh_6_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_440_0 <= mesh_7_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_440_1 <= mesh_7_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_441_0 <= mesh_8_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_441_1 <= mesh_8_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_442_0 <= mesh_9_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_442_1 <= mesh_9_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_443_0 <= mesh_10_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_443_1 <= mesh_10_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_444_0 <= mesh_11_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_444_1 <= mesh_11_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_445_0 <= mesh_12_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_445_1 <= mesh_12_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_446_0 <= mesh_13_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_446_1 <= mesh_13_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_447_0 <= mesh_14_11_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_447_1 <= mesh_14_11_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_448_0 <= io_in_valid_12_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_448_1 <= io_in_valid_12_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_449_0 <= mesh_0_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_449_1 <= mesh_0_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_450_0 <= mesh_1_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_450_1 <= mesh_1_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_451_0 <= mesh_2_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_451_1 <= mesh_2_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_452_0 <= mesh_3_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_452_1 <= mesh_3_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_453_0 <= mesh_4_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_453_1 <= mesh_4_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_454_0 <= mesh_5_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_454_1 <= mesh_5_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_455_0 <= mesh_6_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_455_1 <= mesh_6_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_456_0 <= mesh_7_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_456_1 <= mesh_7_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_457_0 <= mesh_8_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_457_1 <= mesh_8_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_458_0 <= mesh_9_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_458_1 <= mesh_9_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_459_0 <= mesh_10_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_459_1 <= mesh_10_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_460_0 <= mesh_11_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_460_1 <= mesh_11_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_461_0 <= mesh_12_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_461_1 <= mesh_12_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_462_0 <= mesh_13_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_462_1 <= mesh_13_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_463_0 <= mesh_14_12_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_463_1 <= mesh_14_12_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_464_0 <= io_in_valid_13_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_464_1 <= io_in_valid_13_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_465_0 <= mesh_0_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_465_1 <= mesh_0_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_466_0 <= mesh_1_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_466_1 <= mesh_1_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_467_0 <= mesh_2_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_467_1 <= mesh_2_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_468_0 <= mesh_3_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_468_1 <= mesh_3_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_469_0 <= mesh_4_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_469_1 <= mesh_4_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_470_0 <= mesh_5_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_470_1 <= mesh_5_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_471_0 <= mesh_6_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_471_1 <= mesh_6_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_472_0 <= mesh_7_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_472_1 <= mesh_7_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_473_0 <= mesh_8_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_473_1 <= mesh_8_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_474_0 <= mesh_9_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_474_1 <= mesh_9_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_475_0 <= mesh_10_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_475_1 <= mesh_10_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_476_0 <= mesh_11_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_476_1 <= mesh_11_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_477_0 <= mesh_12_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_477_1 <= mesh_12_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_478_0 <= mesh_13_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_478_1 <= mesh_13_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_479_0 <= mesh_14_13_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_479_1 <= mesh_14_13_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_480_0 <= io_in_valid_14_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_480_1 <= io_in_valid_14_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_481_0 <= mesh_0_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_481_1 <= mesh_0_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_482_0 <= mesh_1_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_482_1 <= mesh_1_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_483_0 <= mesh_2_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_483_1 <= mesh_2_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_484_0 <= mesh_3_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_484_1 <= mesh_3_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_485_0 <= mesh_4_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_485_1 <= mesh_4_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_486_0 <= mesh_5_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_486_1 <= mesh_5_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_487_0 <= mesh_6_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_487_1 <= mesh_6_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_488_0 <= mesh_7_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_488_1 <= mesh_7_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_489_0 <= mesh_8_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_489_1 <= mesh_8_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_490_0 <= mesh_9_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_490_1 <= mesh_9_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_491_0 <= mesh_10_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_491_1 <= mesh_10_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_492_0 <= mesh_11_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_492_1 <= mesh_11_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_493_0 <= mesh_12_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_493_1 <= mesh_12_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_494_0 <= mesh_13_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_494_1 <= mesh_13_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_495_0 <= mesh_14_14_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_495_1 <= mesh_14_14_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_496_0 <= io_in_valid_15_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_496_1 <= io_in_valid_15_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_497_0 <= mesh_0_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_497_1 <= mesh_0_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_498_0 <= mesh_1_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_498_1 <= mesh_1_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_499_0 <= mesh_2_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_499_1 <= mesh_2_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_500_0 <= mesh_3_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_500_1 <= mesh_3_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_501_0 <= mesh_4_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_501_1 <= mesh_4_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_502_0 <= mesh_5_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_502_1 <= mesh_5_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_503_0 <= mesh_6_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_503_1 <= mesh_6_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_504_0 <= mesh_7_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_504_1 <= mesh_7_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_505_0 <= mesh_8_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_505_1 <= mesh_8_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_506_0 <= mesh_9_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_506_1 <= mesh_9_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_507_0 <= mesh_10_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_507_1 <= mesh_10_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_508_0 <= mesh_11_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_508_1 <= mesh_11_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_509_0 <= mesh_12_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_509_1 <= mesh_12_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_510_0 <= mesh_13_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_510_1 <= mesh_13_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_511_0 <= mesh_14_15_io_out_valid_0; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_511_1 <= mesh_14_15_io_out_valid_1; // @[src/main/scala/gemmini/Mesh.scala 94:{42,42,42}]
    r_512_0 <= io_in_id_0_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_512_1 <= io_in_id_0_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_513_0 <= mesh_0_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_513_1 <= mesh_0_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_514_0 <= mesh_1_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_514_1 <= mesh_1_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_515_0 <= mesh_2_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_515_1 <= mesh_2_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_516_0 <= mesh_3_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_516_1 <= mesh_3_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_517_0 <= mesh_4_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_517_1 <= mesh_4_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_518_0 <= mesh_5_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_518_1 <= mesh_5_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_519_0 <= mesh_6_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_519_1 <= mesh_6_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_520_0 <= mesh_7_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_520_1 <= mesh_7_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_521_0 <= mesh_8_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_521_1 <= mesh_8_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_522_0 <= mesh_9_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_522_1 <= mesh_9_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_523_0 <= mesh_10_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_523_1 <= mesh_10_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_524_0 <= mesh_11_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_524_1 <= mesh_11_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_525_0 <= mesh_12_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_525_1 <= mesh_12_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_526_0 <= mesh_13_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_526_1 <= mesh_13_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_527_0 <= mesh_14_0_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_527_1 <= mesh_14_0_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_528_0 <= io_in_id_1_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_528_1 <= io_in_id_1_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_529_0 <= mesh_0_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_529_1 <= mesh_0_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_530_0 <= mesh_1_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_530_1 <= mesh_1_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_531_0 <= mesh_2_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_531_1 <= mesh_2_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_532_0 <= mesh_3_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_532_1 <= mesh_3_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_533_0 <= mesh_4_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_533_1 <= mesh_4_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_534_0 <= mesh_5_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_534_1 <= mesh_5_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_535_0 <= mesh_6_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_535_1 <= mesh_6_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_536_0 <= mesh_7_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_536_1 <= mesh_7_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_537_0 <= mesh_8_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_537_1 <= mesh_8_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_538_0 <= mesh_9_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_538_1 <= mesh_9_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_539_0 <= mesh_10_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_539_1 <= mesh_10_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_540_0 <= mesh_11_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_540_1 <= mesh_11_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_541_0 <= mesh_12_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_541_1 <= mesh_12_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_542_0 <= mesh_13_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_542_1 <= mesh_13_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_543_0 <= mesh_14_1_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_543_1 <= mesh_14_1_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_544_0 <= io_in_id_2_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_544_1 <= io_in_id_2_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_545_0 <= mesh_0_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_545_1 <= mesh_0_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_546_0 <= mesh_1_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_546_1 <= mesh_1_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_547_0 <= mesh_2_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_547_1 <= mesh_2_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_548_0 <= mesh_3_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_548_1 <= mesh_3_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_549_0 <= mesh_4_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_549_1 <= mesh_4_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_550_0 <= mesh_5_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_550_1 <= mesh_5_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_551_0 <= mesh_6_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_551_1 <= mesh_6_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_552_0 <= mesh_7_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_552_1 <= mesh_7_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_553_0 <= mesh_8_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_553_1 <= mesh_8_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_554_0 <= mesh_9_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_554_1 <= mesh_9_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_555_0 <= mesh_10_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_555_1 <= mesh_10_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_556_0 <= mesh_11_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_556_1 <= mesh_11_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_557_0 <= mesh_12_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_557_1 <= mesh_12_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_558_0 <= mesh_13_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_558_1 <= mesh_13_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_559_0 <= mesh_14_2_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_559_1 <= mesh_14_2_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_560_0 <= io_in_id_3_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_560_1 <= io_in_id_3_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_561_0 <= mesh_0_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_561_1 <= mesh_0_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_562_0 <= mesh_1_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_562_1 <= mesh_1_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_563_0 <= mesh_2_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_563_1 <= mesh_2_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_564_0 <= mesh_3_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_564_1 <= mesh_3_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_565_0 <= mesh_4_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_565_1 <= mesh_4_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_566_0 <= mesh_5_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_566_1 <= mesh_5_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_567_0 <= mesh_6_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_567_1 <= mesh_6_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_568_0 <= mesh_7_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_568_1 <= mesh_7_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_569_0 <= mesh_8_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_569_1 <= mesh_8_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_570_0 <= mesh_9_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_570_1 <= mesh_9_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_571_0 <= mesh_10_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_571_1 <= mesh_10_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_572_0 <= mesh_11_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_572_1 <= mesh_11_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_573_0 <= mesh_12_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_573_1 <= mesh_12_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_574_0 <= mesh_13_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_574_1 <= mesh_13_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_575_0 <= mesh_14_3_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_575_1 <= mesh_14_3_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_576_0 <= io_in_id_4_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_576_1 <= io_in_id_4_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_577_0 <= mesh_0_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_577_1 <= mesh_0_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_578_0 <= mesh_1_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_578_1 <= mesh_1_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_579_0 <= mesh_2_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_579_1 <= mesh_2_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_580_0 <= mesh_3_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_580_1 <= mesh_3_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_581_0 <= mesh_4_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_581_1 <= mesh_4_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_582_0 <= mesh_5_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_582_1 <= mesh_5_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_583_0 <= mesh_6_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_583_1 <= mesh_6_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_584_0 <= mesh_7_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_584_1 <= mesh_7_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_585_0 <= mesh_8_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_585_1 <= mesh_8_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_586_0 <= mesh_9_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_586_1 <= mesh_9_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_587_0 <= mesh_10_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_587_1 <= mesh_10_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_588_0 <= mesh_11_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_588_1 <= mesh_11_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_589_0 <= mesh_12_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_589_1 <= mesh_12_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_590_0 <= mesh_13_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_590_1 <= mesh_13_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_591_0 <= mesh_14_4_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_591_1 <= mesh_14_4_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_592_0 <= io_in_id_5_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_592_1 <= io_in_id_5_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_593_0 <= mesh_0_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_593_1 <= mesh_0_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_594_0 <= mesh_1_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_594_1 <= mesh_1_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_595_0 <= mesh_2_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_595_1 <= mesh_2_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_596_0 <= mesh_3_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_596_1 <= mesh_3_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_597_0 <= mesh_4_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_597_1 <= mesh_4_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_598_0 <= mesh_5_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_598_1 <= mesh_5_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_599_0 <= mesh_6_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_599_1 <= mesh_6_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_600_0 <= mesh_7_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_600_1 <= mesh_7_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_601_0 <= mesh_8_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_601_1 <= mesh_8_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_602_0 <= mesh_9_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_602_1 <= mesh_9_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_603_0 <= mesh_10_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_603_1 <= mesh_10_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_604_0 <= mesh_11_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_604_1 <= mesh_11_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_605_0 <= mesh_12_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_605_1 <= mesh_12_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_606_0 <= mesh_13_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_606_1 <= mesh_13_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_607_0 <= mesh_14_5_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_607_1 <= mesh_14_5_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_608_0 <= io_in_id_6_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_608_1 <= io_in_id_6_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_609_0 <= mesh_0_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_609_1 <= mesh_0_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_610_0 <= mesh_1_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_610_1 <= mesh_1_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_611_0 <= mesh_2_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_611_1 <= mesh_2_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_612_0 <= mesh_3_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_612_1 <= mesh_3_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_613_0 <= mesh_4_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_613_1 <= mesh_4_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_614_0 <= mesh_5_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_614_1 <= mesh_5_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_615_0 <= mesh_6_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_615_1 <= mesh_6_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_616_0 <= mesh_7_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_616_1 <= mesh_7_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_617_0 <= mesh_8_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_617_1 <= mesh_8_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_618_0 <= mesh_9_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_618_1 <= mesh_9_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_619_0 <= mesh_10_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_619_1 <= mesh_10_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_620_0 <= mesh_11_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_620_1 <= mesh_11_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_621_0 <= mesh_12_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_621_1 <= mesh_12_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_622_0 <= mesh_13_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_622_1 <= mesh_13_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_623_0 <= mesh_14_6_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_623_1 <= mesh_14_6_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_624_0 <= io_in_id_7_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_624_1 <= io_in_id_7_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_625_0 <= mesh_0_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_625_1 <= mesh_0_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_626_0 <= mesh_1_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_626_1 <= mesh_1_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_627_0 <= mesh_2_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_627_1 <= mesh_2_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_628_0 <= mesh_3_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_628_1 <= mesh_3_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_629_0 <= mesh_4_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_629_1 <= mesh_4_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_630_0 <= mesh_5_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_630_1 <= mesh_5_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_631_0 <= mesh_6_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_631_1 <= mesh_6_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_632_0 <= mesh_7_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_632_1 <= mesh_7_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_633_0 <= mesh_8_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_633_1 <= mesh_8_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_634_0 <= mesh_9_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_634_1 <= mesh_9_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_635_0 <= mesh_10_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_635_1 <= mesh_10_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_636_0 <= mesh_11_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_636_1 <= mesh_11_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_637_0 <= mesh_12_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_637_1 <= mesh_12_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_638_0 <= mesh_13_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_638_1 <= mesh_13_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_639_0 <= mesh_14_7_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_639_1 <= mesh_14_7_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_640_0 <= io_in_id_8_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_640_1 <= io_in_id_8_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_641_0 <= mesh_0_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_641_1 <= mesh_0_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_642_0 <= mesh_1_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_642_1 <= mesh_1_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_643_0 <= mesh_2_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_643_1 <= mesh_2_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_644_0 <= mesh_3_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_644_1 <= mesh_3_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_645_0 <= mesh_4_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_645_1 <= mesh_4_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_646_0 <= mesh_5_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_646_1 <= mesh_5_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_647_0 <= mesh_6_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_647_1 <= mesh_6_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_648_0 <= mesh_7_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_648_1 <= mesh_7_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_649_0 <= mesh_8_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_649_1 <= mesh_8_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_650_0 <= mesh_9_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_650_1 <= mesh_9_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_651_0 <= mesh_10_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_651_1 <= mesh_10_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_652_0 <= mesh_11_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_652_1 <= mesh_11_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_653_0 <= mesh_12_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_653_1 <= mesh_12_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_654_0 <= mesh_13_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_654_1 <= mesh_13_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_655_0 <= mesh_14_8_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_655_1 <= mesh_14_8_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_656_0 <= io_in_id_9_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_656_1 <= io_in_id_9_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_657_0 <= mesh_0_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_657_1 <= mesh_0_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_658_0 <= mesh_1_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_658_1 <= mesh_1_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_659_0 <= mesh_2_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_659_1 <= mesh_2_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_660_0 <= mesh_3_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_660_1 <= mesh_3_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_661_0 <= mesh_4_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_661_1 <= mesh_4_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_662_0 <= mesh_5_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_662_1 <= mesh_5_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_663_0 <= mesh_6_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_663_1 <= mesh_6_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_664_0 <= mesh_7_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_664_1 <= mesh_7_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_665_0 <= mesh_8_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_665_1 <= mesh_8_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_666_0 <= mesh_9_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_666_1 <= mesh_9_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_667_0 <= mesh_10_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_667_1 <= mesh_10_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_668_0 <= mesh_11_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_668_1 <= mesh_11_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_669_0 <= mesh_12_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_669_1 <= mesh_12_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_670_0 <= mesh_13_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_670_1 <= mesh_13_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_671_0 <= mesh_14_9_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_671_1 <= mesh_14_9_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_672_0 <= io_in_id_10_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_672_1 <= io_in_id_10_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_673_0 <= mesh_0_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_673_1 <= mesh_0_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_674_0 <= mesh_1_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_674_1 <= mesh_1_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_675_0 <= mesh_2_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_675_1 <= mesh_2_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_676_0 <= mesh_3_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_676_1 <= mesh_3_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_677_0 <= mesh_4_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_677_1 <= mesh_4_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_678_0 <= mesh_5_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_678_1 <= mesh_5_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_679_0 <= mesh_6_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_679_1 <= mesh_6_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_680_0 <= mesh_7_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_680_1 <= mesh_7_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_681_0 <= mesh_8_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_681_1 <= mesh_8_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_682_0 <= mesh_9_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_682_1 <= mesh_9_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_683_0 <= mesh_10_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_683_1 <= mesh_10_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_684_0 <= mesh_11_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_684_1 <= mesh_11_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_685_0 <= mesh_12_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_685_1 <= mesh_12_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_686_0 <= mesh_13_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_686_1 <= mesh_13_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_687_0 <= mesh_14_10_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_687_1 <= mesh_14_10_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_688_0 <= io_in_id_11_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_688_1 <= io_in_id_11_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_689_0 <= mesh_0_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_689_1 <= mesh_0_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_690_0 <= mesh_1_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_690_1 <= mesh_1_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_691_0 <= mesh_2_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_691_1 <= mesh_2_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_692_0 <= mesh_3_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_692_1 <= mesh_3_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_693_0 <= mesh_4_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_693_1 <= mesh_4_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_694_0 <= mesh_5_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_694_1 <= mesh_5_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_695_0 <= mesh_6_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_695_1 <= mesh_6_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_696_0 <= mesh_7_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_696_1 <= mesh_7_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_697_0 <= mesh_8_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_697_1 <= mesh_8_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_698_0 <= mesh_9_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_698_1 <= mesh_9_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_699_0 <= mesh_10_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_699_1 <= mesh_10_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_700_0 <= mesh_11_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_700_1 <= mesh_11_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_701_0 <= mesh_12_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_701_1 <= mesh_12_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_702_0 <= mesh_13_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_702_1 <= mesh_13_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_703_0 <= mesh_14_11_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_703_1 <= mesh_14_11_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_704_0 <= io_in_id_12_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_704_1 <= io_in_id_12_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_705_0 <= mesh_0_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_705_1 <= mesh_0_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_706_0 <= mesh_1_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_706_1 <= mesh_1_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_707_0 <= mesh_2_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_707_1 <= mesh_2_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_708_0 <= mesh_3_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_708_1 <= mesh_3_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_709_0 <= mesh_4_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_709_1 <= mesh_4_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_710_0 <= mesh_5_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_710_1 <= mesh_5_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_711_0 <= mesh_6_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_711_1 <= mesh_6_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_712_0 <= mesh_7_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_712_1 <= mesh_7_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_713_0 <= mesh_8_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_713_1 <= mesh_8_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_714_0 <= mesh_9_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_714_1 <= mesh_9_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_715_0 <= mesh_10_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_715_1 <= mesh_10_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_716_0 <= mesh_11_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_716_1 <= mesh_11_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_717_0 <= mesh_12_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_717_1 <= mesh_12_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_718_0 <= mesh_13_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_718_1 <= mesh_13_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_719_0 <= mesh_14_12_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_719_1 <= mesh_14_12_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_720_0 <= io_in_id_13_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_720_1 <= io_in_id_13_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_721_0 <= mesh_0_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_721_1 <= mesh_0_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_722_0 <= mesh_1_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_722_1 <= mesh_1_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_723_0 <= mesh_2_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_723_1 <= mesh_2_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_724_0 <= mesh_3_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_724_1 <= mesh_3_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_725_0 <= mesh_4_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_725_1 <= mesh_4_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_726_0 <= mesh_5_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_726_1 <= mesh_5_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_727_0 <= mesh_6_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_727_1 <= mesh_6_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_728_0 <= mesh_7_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_728_1 <= mesh_7_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_729_0 <= mesh_8_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_729_1 <= mesh_8_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_730_0 <= mesh_9_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_730_1 <= mesh_9_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_731_0 <= mesh_10_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_731_1 <= mesh_10_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_732_0 <= mesh_11_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_732_1 <= mesh_11_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_733_0 <= mesh_12_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_733_1 <= mesh_12_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_734_0 <= mesh_13_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_734_1 <= mesh_13_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_735_0 <= mesh_14_13_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_735_1 <= mesh_14_13_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_736_0 <= io_in_id_14_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_736_1 <= io_in_id_14_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_737_0 <= mesh_0_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_737_1 <= mesh_0_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_738_0 <= mesh_1_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_738_1 <= mesh_1_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_739_0 <= mesh_2_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_739_1 <= mesh_2_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_740_0 <= mesh_3_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_740_1 <= mesh_3_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_741_0 <= mesh_4_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_741_1 <= mesh_4_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_742_0 <= mesh_5_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_742_1 <= mesh_5_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_743_0 <= mesh_6_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_743_1 <= mesh_6_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_744_0 <= mesh_7_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_744_1 <= mesh_7_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_745_0 <= mesh_8_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_745_1 <= mesh_8_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_746_0 <= mesh_9_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_746_1 <= mesh_9_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_747_0 <= mesh_10_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_747_1 <= mesh_10_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_748_0 <= mesh_11_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_748_1 <= mesh_11_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_749_0 <= mesh_12_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_749_1 <= mesh_12_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_750_0 <= mesh_13_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_750_1 <= mesh_13_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_751_0 <= mesh_14_14_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_751_1 <= mesh_14_14_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_752_0 <= io_in_id_15_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_752_1 <= io_in_id_15_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_753_0 <= mesh_0_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_753_1 <= mesh_0_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_754_0 <= mesh_1_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_754_1 <= mesh_1_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_755_0 <= mesh_2_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_755_1 <= mesh_2_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_756_0 <= mesh_3_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_756_1 <= mesh_3_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_757_0 <= mesh_4_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_757_1 <= mesh_4_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_758_0 <= mesh_5_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_758_1 <= mesh_5_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_759_0 <= mesh_6_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_759_1 <= mesh_6_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_760_0 <= mesh_7_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_760_1 <= mesh_7_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_761_0 <= mesh_8_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_761_1 <= mesh_8_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_762_0 <= mesh_9_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_762_1 <= mesh_9_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_763_0 <= mesh_10_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_763_1 <= mesh_10_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_764_0 <= mesh_11_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_764_1 <= mesh_11_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_765_0 <= mesh_12_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_765_1 <= mesh_12_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_766_0 <= mesh_13_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_766_1 <= mesh_13_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_767_0 <= mesh_14_15_io_out_id_0; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_767_1 <= mesh_14_15_io_out_id_1; // @[src/main/scala/gemmini/Mesh.scala 103:{39,39,39}]
    r_768_0 <= io_in_last_0_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_768_1 <= io_in_last_0_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_769_0 <= mesh_0_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_769_1 <= mesh_0_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_770_0 <= mesh_1_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_770_1 <= mesh_1_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_771_0 <= mesh_2_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_771_1 <= mesh_2_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_772_0 <= mesh_3_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_772_1 <= mesh_3_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_773_0 <= mesh_4_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_773_1 <= mesh_4_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_774_0 <= mesh_5_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_774_1 <= mesh_5_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_775_0 <= mesh_6_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_775_1 <= mesh_6_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_776_0 <= mesh_7_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_776_1 <= mesh_7_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_777_0 <= mesh_8_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_777_1 <= mesh_8_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_778_0 <= mesh_9_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_778_1 <= mesh_9_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_779_0 <= mesh_10_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_779_1 <= mesh_10_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_780_0 <= mesh_11_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_780_1 <= mesh_11_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_781_0 <= mesh_12_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_781_1 <= mesh_12_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_782_0 <= mesh_13_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_782_1 <= mesh_13_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_783_0 <= mesh_14_0_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_783_1 <= mesh_14_0_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_784_0 <= io_in_last_1_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_784_1 <= io_in_last_1_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_785_0 <= mesh_0_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_785_1 <= mesh_0_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_786_0 <= mesh_1_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_786_1 <= mesh_1_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_787_0 <= mesh_2_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_787_1 <= mesh_2_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_788_0 <= mesh_3_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_788_1 <= mesh_3_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_789_0 <= mesh_4_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_789_1 <= mesh_4_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_790_0 <= mesh_5_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_790_1 <= mesh_5_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_791_0 <= mesh_6_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_791_1 <= mesh_6_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_792_0 <= mesh_7_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_792_1 <= mesh_7_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_793_0 <= mesh_8_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_793_1 <= mesh_8_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_794_0 <= mesh_9_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_794_1 <= mesh_9_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_795_0 <= mesh_10_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_795_1 <= mesh_10_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_796_0 <= mesh_11_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_796_1 <= mesh_11_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_797_0 <= mesh_12_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_797_1 <= mesh_12_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_798_0 <= mesh_13_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_798_1 <= mesh_13_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_799_0 <= mesh_14_1_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_799_1 <= mesh_14_1_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_800_0 <= io_in_last_2_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_800_1 <= io_in_last_2_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_801_0 <= mesh_0_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_801_1 <= mesh_0_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_802_0 <= mesh_1_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_802_1 <= mesh_1_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_803_0 <= mesh_2_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_803_1 <= mesh_2_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_804_0 <= mesh_3_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_804_1 <= mesh_3_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_805_0 <= mesh_4_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_805_1 <= mesh_4_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_806_0 <= mesh_5_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_806_1 <= mesh_5_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_807_0 <= mesh_6_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_807_1 <= mesh_6_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_808_0 <= mesh_7_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_808_1 <= mesh_7_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_809_0 <= mesh_8_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_809_1 <= mesh_8_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_810_0 <= mesh_9_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_810_1 <= mesh_9_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_811_0 <= mesh_10_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_811_1 <= mesh_10_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_812_0 <= mesh_11_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_812_1 <= mesh_11_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_813_0 <= mesh_12_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_813_1 <= mesh_12_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_814_0 <= mesh_13_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_814_1 <= mesh_13_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_815_0 <= mesh_14_2_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_815_1 <= mesh_14_2_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_816_0 <= io_in_last_3_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_816_1 <= io_in_last_3_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_817_0 <= mesh_0_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_817_1 <= mesh_0_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_818_0 <= mesh_1_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_818_1 <= mesh_1_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_819_0 <= mesh_2_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_819_1 <= mesh_2_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_820_0 <= mesh_3_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_820_1 <= mesh_3_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_821_0 <= mesh_4_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_821_1 <= mesh_4_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_822_0 <= mesh_5_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_822_1 <= mesh_5_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_823_0 <= mesh_6_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_823_1 <= mesh_6_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_824_0 <= mesh_7_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_824_1 <= mesh_7_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_825_0 <= mesh_8_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_825_1 <= mesh_8_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_826_0 <= mesh_9_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_826_1 <= mesh_9_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_827_0 <= mesh_10_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_827_1 <= mesh_10_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_828_0 <= mesh_11_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_828_1 <= mesh_11_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_829_0 <= mesh_12_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_829_1 <= mesh_12_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_830_0 <= mesh_13_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_830_1 <= mesh_13_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_831_0 <= mesh_14_3_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_831_1 <= mesh_14_3_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_832_0 <= io_in_last_4_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_832_1 <= io_in_last_4_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_833_0 <= mesh_0_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_833_1 <= mesh_0_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_834_0 <= mesh_1_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_834_1 <= mesh_1_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_835_0 <= mesh_2_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_835_1 <= mesh_2_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_836_0 <= mesh_3_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_836_1 <= mesh_3_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_837_0 <= mesh_4_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_837_1 <= mesh_4_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_838_0 <= mesh_5_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_838_1 <= mesh_5_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_839_0 <= mesh_6_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_839_1 <= mesh_6_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_840_0 <= mesh_7_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_840_1 <= mesh_7_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_841_0 <= mesh_8_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_841_1 <= mesh_8_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_842_0 <= mesh_9_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_842_1 <= mesh_9_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_843_0 <= mesh_10_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_843_1 <= mesh_10_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_844_0 <= mesh_11_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_844_1 <= mesh_11_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_845_0 <= mesh_12_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_845_1 <= mesh_12_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_846_0 <= mesh_13_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_846_1 <= mesh_13_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_847_0 <= mesh_14_4_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_847_1 <= mesh_14_4_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_848_0 <= io_in_last_5_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_848_1 <= io_in_last_5_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_849_0 <= mesh_0_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_849_1 <= mesh_0_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_850_0 <= mesh_1_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_850_1 <= mesh_1_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_851_0 <= mesh_2_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_851_1 <= mesh_2_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_852_0 <= mesh_3_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_852_1 <= mesh_3_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_853_0 <= mesh_4_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_853_1 <= mesh_4_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_854_0 <= mesh_5_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_854_1 <= mesh_5_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_855_0 <= mesh_6_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_855_1 <= mesh_6_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_856_0 <= mesh_7_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_856_1 <= mesh_7_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_857_0 <= mesh_8_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_857_1 <= mesh_8_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_858_0 <= mesh_9_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_858_1 <= mesh_9_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_859_0 <= mesh_10_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_859_1 <= mesh_10_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_860_0 <= mesh_11_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_860_1 <= mesh_11_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_861_0 <= mesh_12_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_861_1 <= mesh_12_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_862_0 <= mesh_13_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_862_1 <= mesh_13_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_863_0 <= mesh_14_5_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_863_1 <= mesh_14_5_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_864_0 <= io_in_last_6_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_864_1 <= io_in_last_6_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_865_0 <= mesh_0_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_865_1 <= mesh_0_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_866_0 <= mesh_1_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_866_1 <= mesh_1_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_867_0 <= mesh_2_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_867_1 <= mesh_2_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_868_0 <= mesh_3_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_868_1 <= mesh_3_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_869_0 <= mesh_4_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_869_1 <= mesh_4_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_870_0 <= mesh_5_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_870_1 <= mesh_5_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_871_0 <= mesh_6_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_871_1 <= mesh_6_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_872_0 <= mesh_7_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_872_1 <= mesh_7_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_873_0 <= mesh_8_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_873_1 <= mesh_8_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_874_0 <= mesh_9_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_874_1 <= mesh_9_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_875_0 <= mesh_10_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_875_1 <= mesh_10_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_876_0 <= mesh_11_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_876_1 <= mesh_11_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_877_0 <= mesh_12_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_877_1 <= mesh_12_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_878_0 <= mesh_13_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_878_1 <= mesh_13_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_879_0 <= mesh_14_6_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_879_1 <= mesh_14_6_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_880_0 <= io_in_last_7_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_880_1 <= io_in_last_7_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_881_0 <= mesh_0_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_881_1 <= mesh_0_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_882_0 <= mesh_1_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_882_1 <= mesh_1_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_883_0 <= mesh_2_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_883_1 <= mesh_2_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_884_0 <= mesh_3_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_884_1 <= mesh_3_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_885_0 <= mesh_4_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_885_1 <= mesh_4_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_886_0 <= mesh_5_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_886_1 <= mesh_5_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_887_0 <= mesh_6_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_887_1 <= mesh_6_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_888_0 <= mesh_7_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_888_1 <= mesh_7_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_889_0 <= mesh_8_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_889_1 <= mesh_8_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_890_0 <= mesh_9_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_890_1 <= mesh_9_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_891_0 <= mesh_10_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_891_1 <= mesh_10_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_892_0 <= mesh_11_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_892_1 <= mesh_11_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_893_0 <= mesh_12_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_893_1 <= mesh_12_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_894_0 <= mesh_13_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_894_1 <= mesh_13_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_895_0 <= mesh_14_7_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_895_1 <= mesh_14_7_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_896_0 <= io_in_last_8_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_896_1 <= io_in_last_8_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_897_0 <= mesh_0_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_897_1 <= mesh_0_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_898_0 <= mesh_1_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_898_1 <= mesh_1_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_899_0 <= mesh_2_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_899_1 <= mesh_2_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_900_0 <= mesh_3_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_900_1 <= mesh_3_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_901_0 <= mesh_4_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_901_1 <= mesh_4_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_902_0 <= mesh_5_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_902_1 <= mesh_5_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_903_0 <= mesh_6_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_903_1 <= mesh_6_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_904_0 <= mesh_7_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_904_1 <= mesh_7_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_905_0 <= mesh_8_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_905_1 <= mesh_8_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_906_0 <= mesh_9_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_906_1 <= mesh_9_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_907_0 <= mesh_10_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_907_1 <= mesh_10_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_908_0 <= mesh_11_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_908_1 <= mesh_11_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_909_0 <= mesh_12_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_909_1 <= mesh_12_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_910_0 <= mesh_13_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_910_1 <= mesh_13_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_911_0 <= mesh_14_8_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_911_1 <= mesh_14_8_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_912_0 <= io_in_last_9_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_912_1 <= io_in_last_9_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_913_0 <= mesh_0_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_913_1 <= mesh_0_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_914_0 <= mesh_1_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_914_1 <= mesh_1_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_915_0 <= mesh_2_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_915_1 <= mesh_2_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_916_0 <= mesh_3_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_916_1 <= mesh_3_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_917_0 <= mesh_4_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_917_1 <= mesh_4_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_918_0 <= mesh_5_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_918_1 <= mesh_5_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_919_0 <= mesh_6_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_919_1 <= mesh_6_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_920_0 <= mesh_7_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_920_1 <= mesh_7_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_921_0 <= mesh_8_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_921_1 <= mesh_8_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_922_0 <= mesh_9_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_922_1 <= mesh_9_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_923_0 <= mesh_10_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_923_1 <= mesh_10_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_924_0 <= mesh_11_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_924_1 <= mesh_11_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_925_0 <= mesh_12_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_925_1 <= mesh_12_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_926_0 <= mesh_13_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_926_1 <= mesh_13_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_927_0 <= mesh_14_9_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_927_1 <= mesh_14_9_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_928_0 <= io_in_last_10_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_928_1 <= io_in_last_10_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_929_0 <= mesh_0_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_929_1 <= mesh_0_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_930_0 <= mesh_1_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_930_1 <= mesh_1_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_931_0 <= mesh_2_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_931_1 <= mesh_2_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_932_0 <= mesh_3_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_932_1 <= mesh_3_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_933_0 <= mesh_4_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_933_1 <= mesh_4_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_934_0 <= mesh_5_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_934_1 <= mesh_5_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_935_0 <= mesh_6_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_935_1 <= mesh_6_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_936_0 <= mesh_7_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_936_1 <= mesh_7_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_937_0 <= mesh_8_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_937_1 <= mesh_8_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_938_0 <= mesh_9_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_938_1 <= mesh_9_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_939_0 <= mesh_10_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_939_1 <= mesh_10_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_940_0 <= mesh_11_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_940_1 <= mesh_11_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_941_0 <= mesh_12_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_941_1 <= mesh_12_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_942_0 <= mesh_13_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_942_1 <= mesh_13_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_943_0 <= mesh_14_10_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_943_1 <= mesh_14_10_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_944_0 <= io_in_last_11_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_944_1 <= io_in_last_11_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_945_0 <= mesh_0_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_945_1 <= mesh_0_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_946_0 <= mesh_1_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_946_1 <= mesh_1_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_947_0 <= mesh_2_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_947_1 <= mesh_2_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_948_0 <= mesh_3_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_948_1 <= mesh_3_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_949_0 <= mesh_4_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_949_1 <= mesh_4_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_950_0 <= mesh_5_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_950_1 <= mesh_5_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_951_0 <= mesh_6_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_951_1 <= mesh_6_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_952_0 <= mesh_7_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_952_1 <= mesh_7_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_953_0 <= mesh_8_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_953_1 <= mesh_8_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_954_0 <= mesh_9_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_954_1 <= mesh_9_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_955_0 <= mesh_10_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_955_1 <= mesh_10_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_956_0 <= mesh_11_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_956_1 <= mesh_11_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_957_0 <= mesh_12_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_957_1 <= mesh_12_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_958_0 <= mesh_13_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_958_1 <= mesh_13_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_959_0 <= mesh_14_11_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_959_1 <= mesh_14_11_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_960_0 <= io_in_last_12_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_960_1 <= io_in_last_12_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_961_0 <= mesh_0_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_961_1 <= mesh_0_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_962_0 <= mesh_1_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_962_1 <= mesh_1_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_963_0 <= mesh_2_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_963_1 <= mesh_2_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_964_0 <= mesh_3_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_964_1 <= mesh_3_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_965_0 <= mesh_4_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_965_1 <= mesh_4_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_966_0 <= mesh_5_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_966_1 <= mesh_5_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_967_0 <= mesh_6_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_967_1 <= mesh_6_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_968_0 <= mesh_7_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_968_1 <= mesh_7_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_969_0 <= mesh_8_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_969_1 <= mesh_8_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_970_0 <= mesh_9_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_970_1 <= mesh_9_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_971_0 <= mesh_10_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_971_1 <= mesh_10_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_972_0 <= mesh_11_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_972_1 <= mesh_11_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_973_0 <= mesh_12_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_973_1 <= mesh_12_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_974_0 <= mesh_13_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_974_1 <= mesh_13_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_975_0 <= mesh_14_12_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_975_1 <= mesh_14_12_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_976_0 <= io_in_last_13_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_976_1 <= io_in_last_13_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_977_0 <= mesh_0_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_977_1 <= mesh_0_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_978_0 <= mesh_1_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_978_1 <= mesh_1_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_979_0 <= mesh_2_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_979_1 <= mesh_2_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_980_0 <= mesh_3_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_980_1 <= mesh_3_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_981_0 <= mesh_4_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_981_1 <= mesh_4_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_982_0 <= mesh_5_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_982_1 <= mesh_5_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_983_0 <= mesh_6_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_983_1 <= mesh_6_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_984_0 <= mesh_7_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_984_1 <= mesh_7_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_985_0 <= mesh_8_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_985_1 <= mesh_8_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_986_0 <= mesh_9_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_986_1 <= mesh_9_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_987_0 <= mesh_10_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_987_1 <= mesh_10_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_988_0 <= mesh_11_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_988_1 <= mesh_11_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_989_0 <= mesh_12_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_989_1 <= mesh_12_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_990_0 <= mesh_13_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_990_1 <= mesh_13_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_991_0 <= mesh_14_13_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_991_1 <= mesh_14_13_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_992_0 <= io_in_last_14_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_992_1 <= io_in_last_14_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_993_0 <= mesh_0_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_993_1 <= mesh_0_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_994_0 <= mesh_1_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_994_1 <= mesh_1_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_995_0 <= mesh_2_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_995_1 <= mesh_2_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_996_0 <= mesh_3_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_996_1 <= mesh_3_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_997_0 <= mesh_4_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_997_1 <= mesh_4_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_998_0 <= mesh_5_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_998_1 <= mesh_5_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_999_0 <= mesh_6_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_999_1 <= mesh_6_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1000_0 <= mesh_7_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1000_1 <= mesh_7_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1001_0 <= mesh_8_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1001_1 <= mesh_8_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1002_0 <= mesh_9_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1002_1 <= mesh_9_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1003_0 <= mesh_10_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1003_1 <= mesh_10_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1004_0 <= mesh_11_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1004_1 <= mesh_11_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1005_0 <= mesh_12_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1005_1 <= mesh_12_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1006_0 <= mesh_13_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1006_1 <= mesh_13_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1007_0 <= mesh_14_14_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1007_1 <= mesh_14_14_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1008_0 <= io_in_last_15_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1008_1 <= io_in_last_15_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1009_0 <= mesh_0_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1009_1 <= mesh_0_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1010_0 <= mesh_1_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1010_1 <= mesh_1_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1011_0 <= mesh_2_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1011_1 <= mesh_2_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1012_0 <= mesh_3_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1012_1 <= mesh_3_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1013_0 <= mesh_4_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1013_1 <= mesh_4_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1014_0 <= mesh_5_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1014_1 <= mesh_5_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1015_0 <= mesh_6_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1015_1 <= mesh_6_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1016_0 <= mesh_7_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1016_1 <= mesh_7_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1017_0 <= mesh_8_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1017_1 <= mesh_8_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1018_0 <= mesh_9_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1018_1 <= mesh_9_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1019_0 <= mesh_10_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1019_1 <= mesh_10_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1020_0 <= mesh_11_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1020_1 <= mesh_11_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1021_0 <= mesh_12_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1021_1 <= mesh_12_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1022_0 <= mesh_13_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1022_1 <= mesh_13_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1023_0 <= mesh_14_15_io_out_last_0; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
    r_1023_1 <= mesh_14_15_io_out_last_1; // @[src/main/scala/gemmini/Mesh.scala 112:{41,41,41}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r__0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  r__1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  r_1_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  r_1_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  r_2_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  r_2_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_3_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_3_1 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_4_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r_4_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  r_5_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  r_5_1 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_6_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  r_6_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  r_7_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  r_7_1 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  r_8_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  r_8_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  r_9_0 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  r_9_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  r_10_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  r_10_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  r_11_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  r_11_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  r_12_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  r_12_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  r_13_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  r_13_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  r_14_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  r_14_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  r_15_0 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  r_15_1 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  r_16_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  r_16_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  r_17_0 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  r_17_1 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  r_18_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  r_18_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  r_19_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  r_19_1 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  r_20_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  r_20_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  r_21_0 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  r_21_1 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  r_22_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  r_22_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  r_23_0 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  r_23_1 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  r_24_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  r_24_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  r_25_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  r_25_1 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  r_26_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  r_26_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  r_27_0 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  r_27_1 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  r_28_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  r_28_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  r_29_0 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  r_29_1 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  r_30_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  r_30_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  r_31_0 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  r_31_1 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  r_32_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  r_32_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  r_33_0 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  r_33_1 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  r_34_0 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  r_34_1 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  r_35_0 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  r_35_1 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  r_36_0 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  r_36_1 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  r_37_0 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  r_37_1 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  r_38_0 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  r_38_1 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  r_39_0 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  r_39_1 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  r_40_0 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  r_40_1 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  r_41_0 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  r_41_1 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  r_42_0 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  r_42_1 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  r_43_0 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  r_43_1 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  r_44_0 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  r_44_1 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  r_45_0 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  r_45_1 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  r_46_0 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  r_46_1 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  r_47_0 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  r_47_1 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  r_48_0 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  r_48_1 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  r_49_0 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  r_49_1 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  r_50_0 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  r_50_1 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  r_51_0 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  r_51_1 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  r_52_0 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  r_52_1 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  r_53_0 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  r_53_1 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  r_54_0 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  r_54_1 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  r_55_0 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  r_55_1 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  r_56_0 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  r_56_1 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  r_57_0 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  r_57_1 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  r_58_0 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  r_58_1 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  r_59_0 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  r_59_1 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  r_60_0 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  r_60_1 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  r_61_0 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  r_61_1 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  r_62_0 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  r_62_1 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  r_63_0 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  r_63_1 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  r_64_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  r_64_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  r_65_0 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  r_65_1 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  r_66_0 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  r_66_1 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  r_67_0 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  r_67_1 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  r_68_0 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  r_68_1 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  r_69_0 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  r_69_1 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  r_70_0 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  r_70_1 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  r_71_0 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  r_71_1 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  r_72_0 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  r_72_1 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  r_73_0 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  r_73_1 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  r_74_0 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  r_74_1 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  r_75_0 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  r_75_1 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  r_76_0 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  r_76_1 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  r_77_0 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  r_77_1 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  r_78_0 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  r_78_1 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  r_79_0 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  r_79_1 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  r_80_0 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  r_80_1 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  r_81_0 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  r_81_1 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  r_82_0 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  r_82_1 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  r_83_0 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  r_83_1 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  r_84_0 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  r_84_1 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  r_85_0 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  r_85_1 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  r_86_0 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  r_86_1 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  r_87_0 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  r_87_1 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  r_88_0 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  r_88_1 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  r_89_0 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  r_89_1 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  r_90_0 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  r_90_1 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  r_91_0 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  r_91_1 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  r_92_0 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  r_92_1 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  r_93_0 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  r_93_1 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  r_94_0 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  r_94_1 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  r_95_0 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  r_95_1 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  r_96_0 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  r_96_1 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  r_97_0 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  r_97_1 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  r_98_0 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  r_98_1 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  r_99_0 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  r_99_1 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  r_100_0 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  r_100_1 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  r_101_0 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  r_101_1 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  r_102_0 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  r_102_1 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  r_103_0 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  r_103_1 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  r_104_0 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  r_104_1 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  r_105_0 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  r_105_1 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  r_106_0 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  r_106_1 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  r_107_0 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  r_107_1 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  r_108_0 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  r_108_1 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  r_109_0 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  r_109_1 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  r_110_0 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  r_110_1 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  r_111_0 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  r_111_1 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  r_112_0 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  r_112_1 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  r_113_0 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  r_113_1 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  r_114_0 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  r_114_1 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  r_115_0 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  r_115_1 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  r_116_0 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  r_116_1 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  r_117_0 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  r_117_1 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  r_118_0 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  r_118_1 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  r_119_0 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  r_119_1 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  r_120_0 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  r_120_1 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  r_121_0 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  r_121_1 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  r_122_0 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  r_122_1 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  r_123_0 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  r_123_1 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  r_124_0 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  r_124_1 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  r_125_0 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  r_125_1 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  r_126_0 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  r_126_1 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  r_127_0 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  r_127_1 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  r_128_0 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  r_128_1 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  r_129_0 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  r_129_1 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  r_130_0 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  r_130_1 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  r_131_0 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  r_131_1 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  r_132_0 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  r_132_1 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  r_133_0 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  r_133_1 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  r_134_0 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  r_134_1 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  r_135_0 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  r_135_1 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  r_136_0 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  r_136_1 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  r_137_0 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  r_137_1 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  r_138_0 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  r_138_1 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  r_139_0 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  r_139_1 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  r_140_0 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  r_140_1 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  r_141_0 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  r_141_1 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  r_142_0 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  r_142_1 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  r_143_0 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  r_143_1 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  r_144_0 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  r_144_1 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  r_145_0 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  r_145_1 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  r_146_0 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  r_146_1 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  r_147_0 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  r_147_1 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  r_148_0 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  r_148_1 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  r_149_0 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  r_149_1 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  r_150_0 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  r_150_1 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  r_151_0 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  r_151_1 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  r_152_0 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  r_152_1 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  r_153_0 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  r_153_1 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  r_154_0 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  r_154_1 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  r_155_0 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  r_155_1 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  r_156_0 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  r_156_1 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  r_157_0 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  r_157_1 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  r_158_0 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  r_158_1 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  r_159_0 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  r_159_1 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  r_160_0 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  r_160_1 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  r_161_0 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  r_161_1 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  r_162_0 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  r_162_1 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  r_163_0 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  r_163_1 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  r_164_0 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  r_164_1 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  r_165_0 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  r_165_1 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  r_166_0 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  r_166_1 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  r_167_0 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  r_167_1 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  r_168_0 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  r_168_1 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  r_169_0 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  r_169_1 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  r_170_0 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  r_170_1 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  r_171_0 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  r_171_1 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  r_172_0 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  r_172_1 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  r_173_0 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  r_173_1 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  r_174_0 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  r_174_1 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  r_175_0 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  r_175_1 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  r_176_0 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  r_176_1 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  r_177_0 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  r_177_1 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  r_178_0 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  r_178_1 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  r_179_0 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  r_179_1 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  r_180_0 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  r_180_1 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  r_181_0 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  r_181_1 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  r_182_0 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  r_182_1 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  r_183_0 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  r_183_1 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  r_184_0 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  r_184_1 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  r_185_0 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  r_185_1 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  r_186_0 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  r_186_1 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  r_187_0 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  r_187_1 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  r_188_0 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  r_188_1 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  r_189_0 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  r_189_1 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  r_190_0 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  r_190_1 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  r_191_0 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  r_191_1 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  r_192_0 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  r_192_1 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  r_193_0 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  r_193_1 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  r_194_0 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  r_194_1 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  r_195_0 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  r_195_1 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  r_196_0 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  r_196_1 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  r_197_0 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  r_197_1 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  r_198_0 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  r_198_1 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  r_199_0 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  r_199_1 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  r_200_0 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  r_200_1 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  r_201_0 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  r_201_1 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  r_202_0 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  r_202_1 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  r_203_0 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  r_203_1 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  r_204_0 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  r_204_1 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  r_205_0 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  r_205_1 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  r_206_0 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  r_206_1 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  r_207_0 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  r_207_1 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  r_208_0 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  r_208_1 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  r_209_0 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  r_209_1 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  r_210_0 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  r_210_1 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  r_211_0 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  r_211_1 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  r_212_0 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  r_212_1 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  r_213_0 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  r_213_1 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  r_214_0 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  r_214_1 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  r_215_0 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  r_215_1 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  r_216_0 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  r_216_1 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  r_217_0 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  r_217_1 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  r_218_0 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  r_218_1 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  r_219_0 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  r_219_1 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  r_220_0 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  r_220_1 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  r_221_0 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  r_221_1 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  r_222_0 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  r_222_1 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  r_223_0 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  r_223_1 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  r_224_0 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  r_224_1 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  r_225_0 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  r_225_1 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  r_226_0 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  r_226_1 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  r_227_0 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  r_227_1 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  r_228_0 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  r_228_1 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  r_229_0 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  r_229_1 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  r_230_0 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  r_230_1 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  r_231_0 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  r_231_1 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  r_232_0 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  r_232_1 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  r_233_0 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  r_233_1 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  r_234_0 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  r_234_1 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  r_235_0 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  r_235_1 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  r_236_0 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  r_236_1 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  r_237_0 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  r_237_1 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  r_238_0 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  r_238_1 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  r_239_0 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  r_239_1 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  r_240_0 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  r_240_1 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  r_241_0 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  r_241_1 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  r_242_0 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  r_242_1 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  r_243_0 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  r_243_1 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  r_244_0 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  r_244_1 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  r_245_0 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  r_245_1 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  r_246_0 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  r_246_1 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  r_247_0 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  r_247_1 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  r_248_0 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  r_248_1 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  r_249_0 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  r_249_1 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  r_250_0 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  r_250_1 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  r_251_0 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  r_251_1 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  r_252_0 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  r_252_1 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  r_253_0 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  r_253_1 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  r_254_0 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  r_254_1 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  r_255_0 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  r_255_1 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  pipe_b__0 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  pipe_b__1 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  pipe_b_1_0 = _RAND_514[19:0];
  _RAND_515 = {1{`RANDOM}};
  pipe_b_1_1 = _RAND_515[19:0];
  _RAND_516 = {1{`RANDOM}};
  pipe_b_2_0 = _RAND_516[19:0];
  _RAND_517 = {1{`RANDOM}};
  pipe_b_2_1 = _RAND_517[19:0];
  _RAND_518 = {1{`RANDOM}};
  pipe_b_3_0 = _RAND_518[19:0];
  _RAND_519 = {1{`RANDOM}};
  pipe_b_3_1 = _RAND_519[19:0];
  _RAND_520 = {1{`RANDOM}};
  pipe_b_4_0 = _RAND_520[19:0];
  _RAND_521 = {1{`RANDOM}};
  pipe_b_4_1 = _RAND_521[19:0];
  _RAND_522 = {1{`RANDOM}};
  pipe_b_5_0 = _RAND_522[19:0];
  _RAND_523 = {1{`RANDOM}};
  pipe_b_5_1 = _RAND_523[19:0];
  _RAND_524 = {1{`RANDOM}};
  pipe_b_6_0 = _RAND_524[19:0];
  _RAND_525 = {1{`RANDOM}};
  pipe_b_6_1 = _RAND_525[19:0];
  _RAND_526 = {1{`RANDOM}};
  pipe_b_7_0 = _RAND_526[19:0];
  _RAND_527 = {1{`RANDOM}};
  pipe_b_7_1 = _RAND_527[19:0];
  _RAND_528 = {1{`RANDOM}};
  pipe_b_8_0 = _RAND_528[19:0];
  _RAND_529 = {1{`RANDOM}};
  pipe_b_8_1 = _RAND_529[19:0];
  _RAND_530 = {1{`RANDOM}};
  pipe_b_9_0 = _RAND_530[19:0];
  _RAND_531 = {1{`RANDOM}};
  pipe_b_9_1 = _RAND_531[19:0];
  _RAND_532 = {1{`RANDOM}};
  pipe_b_10_0 = _RAND_532[19:0];
  _RAND_533 = {1{`RANDOM}};
  pipe_b_10_1 = _RAND_533[19:0];
  _RAND_534 = {1{`RANDOM}};
  pipe_b_11_0 = _RAND_534[19:0];
  _RAND_535 = {1{`RANDOM}};
  pipe_b_11_1 = _RAND_535[19:0];
  _RAND_536 = {1{`RANDOM}};
  pipe_b_12_0 = _RAND_536[19:0];
  _RAND_537 = {1{`RANDOM}};
  pipe_b_12_1 = _RAND_537[19:0];
  _RAND_538 = {1{`RANDOM}};
  pipe_b_13_0 = _RAND_538[19:0];
  _RAND_539 = {1{`RANDOM}};
  pipe_b_13_1 = _RAND_539[19:0];
  _RAND_540 = {1{`RANDOM}};
  pipe_b_14_0 = _RAND_540[19:0];
  _RAND_541 = {1{`RANDOM}};
  pipe_b_14_1 = _RAND_541[19:0];
  _RAND_542 = {1{`RANDOM}};
  pipe_b_15_0 = _RAND_542[19:0];
  _RAND_543 = {1{`RANDOM}};
  pipe_b_15_1 = _RAND_543[19:0];
  _RAND_544 = {1{`RANDOM}};
  pipe_b_16_0 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  pipe_b_16_1 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  pipe_b_17_0 = _RAND_546[19:0];
  _RAND_547 = {1{`RANDOM}};
  pipe_b_17_1 = _RAND_547[19:0];
  _RAND_548 = {1{`RANDOM}};
  pipe_b_18_0 = _RAND_548[19:0];
  _RAND_549 = {1{`RANDOM}};
  pipe_b_18_1 = _RAND_549[19:0];
  _RAND_550 = {1{`RANDOM}};
  pipe_b_19_0 = _RAND_550[19:0];
  _RAND_551 = {1{`RANDOM}};
  pipe_b_19_1 = _RAND_551[19:0];
  _RAND_552 = {1{`RANDOM}};
  pipe_b_20_0 = _RAND_552[19:0];
  _RAND_553 = {1{`RANDOM}};
  pipe_b_20_1 = _RAND_553[19:0];
  _RAND_554 = {1{`RANDOM}};
  pipe_b_21_0 = _RAND_554[19:0];
  _RAND_555 = {1{`RANDOM}};
  pipe_b_21_1 = _RAND_555[19:0];
  _RAND_556 = {1{`RANDOM}};
  pipe_b_22_0 = _RAND_556[19:0];
  _RAND_557 = {1{`RANDOM}};
  pipe_b_22_1 = _RAND_557[19:0];
  _RAND_558 = {1{`RANDOM}};
  pipe_b_23_0 = _RAND_558[19:0];
  _RAND_559 = {1{`RANDOM}};
  pipe_b_23_1 = _RAND_559[19:0];
  _RAND_560 = {1{`RANDOM}};
  pipe_b_24_0 = _RAND_560[19:0];
  _RAND_561 = {1{`RANDOM}};
  pipe_b_24_1 = _RAND_561[19:0];
  _RAND_562 = {1{`RANDOM}};
  pipe_b_25_0 = _RAND_562[19:0];
  _RAND_563 = {1{`RANDOM}};
  pipe_b_25_1 = _RAND_563[19:0];
  _RAND_564 = {1{`RANDOM}};
  pipe_b_26_0 = _RAND_564[19:0];
  _RAND_565 = {1{`RANDOM}};
  pipe_b_26_1 = _RAND_565[19:0];
  _RAND_566 = {1{`RANDOM}};
  pipe_b_27_0 = _RAND_566[19:0];
  _RAND_567 = {1{`RANDOM}};
  pipe_b_27_1 = _RAND_567[19:0];
  _RAND_568 = {1{`RANDOM}};
  pipe_b_28_0 = _RAND_568[19:0];
  _RAND_569 = {1{`RANDOM}};
  pipe_b_28_1 = _RAND_569[19:0];
  _RAND_570 = {1{`RANDOM}};
  pipe_b_29_0 = _RAND_570[19:0];
  _RAND_571 = {1{`RANDOM}};
  pipe_b_29_1 = _RAND_571[19:0];
  _RAND_572 = {1{`RANDOM}};
  pipe_b_30_0 = _RAND_572[19:0];
  _RAND_573 = {1{`RANDOM}};
  pipe_b_30_1 = _RAND_573[19:0];
  _RAND_574 = {1{`RANDOM}};
  pipe_b_31_0 = _RAND_574[19:0];
  _RAND_575 = {1{`RANDOM}};
  pipe_b_31_1 = _RAND_575[19:0];
  _RAND_576 = {1{`RANDOM}};
  pipe_b_32_0 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  pipe_b_32_1 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  pipe_b_33_0 = _RAND_578[19:0];
  _RAND_579 = {1{`RANDOM}};
  pipe_b_33_1 = _RAND_579[19:0];
  _RAND_580 = {1{`RANDOM}};
  pipe_b_34_0 = _RAND_580[19:0];
  _RAND_581 = {1{`RANDOM}};
  pipe_b_34_1 = _RAND_581[19:0];
  _RAND_582 = {1{`RANDOM}};
  pipe_b_35_0 = _RAND_582[19:0];
  _RAND_583 = {1{`RANDOM}};
  pipe_b_35_1 = _RAND_583[19:0];
  _RAND_584 = {1{`RANDOM}};
  pipe_b_36_0 = _RAND_584[19:0];
  _RAND_585 = {1{`RANDOM}};
  pipe_b_36_1 = _RAND_585[19:0];
  _RAND_586 = {1{`RANDOM}};
  pipe_b_37_0 = _RAND_586[19:0];
  _RAND_587 = {1{`RANDOM}};
  pipe_b_37_1 = _RAND_587[19:0];
  _RAND_588 = {1{`RANDOM}};
  pipe_b_38_0 = _RAND_588[19:0];
  _RAND_589 = {1{`RANDOM}};
  pipe_b_38_1 = _RAND_589[19:0];
  _RAND_590 = {1{`RANDOM}};
  pipe_b_39_0 = _RAND_590[19:0];
  _RAND_591 = {1{`RANDOM}};
  pipe_b_39_1 = _RAND_591[19:0];
  _RAND_592 = {1{`RANDOM}};
  pipe_b_40_0 = _RAND_592[19:0];
  _RAND_593 = {1{`RANDOM}};
  pipe_b_40_1 = _RAND_593[19:0];
  _RAND_594 = {1{`RANDOM}};
  pipe_b_41_0 = _RAND_594[19:0];
  _RAND_595 = {1{`RANDOM}};
  pipe_b_41_1 = _RAND_595[19:0];
  _RAND_596 = {1{`RANDOM}};
  pipe_b_42_0 = _RAND_596[19:0];
  _RAND_597 = {1{`RANDOM}};
  pipe_b_42_1 = _RAND_597[19:0];
  _RAND_598 = {1{`RANDOM}};
  pipe_b_43_0 = _RAND_598[19:0];
  _RAND_599 = {1{`RANDOM}};
  pipe_b_43_1 = _RAND_599[19:0];
  _RAND_600 = {1{`RANDOM}};
  pipe_b_44_0 = _RAND_600[19:0];
  _RAND_601 = {1{`RANDOM}};
  pipe_b_44_1 = _RAND_601[19:0];
  _RAND_602 = {1{`RANDOM}};
  pipe_b_45_0 = _RAND_602[19:0];
  _RAND_603 = {1{`RANDOM}};
  pipe_b_45_1 = _RAND_603[19:0];
  _RAND_604 = {1{`RANDOM}};
  pipe_b_46_0 = _RAND_604[19:0];
  _RAND_605 = {1{`RANDOM}};
  pipe_b_46_1 = _RAND_605[19:0];
  _RAND_606 = {1{`RANDOM}};
  pipe_b_47_0 = _RAND_606[19:0];
  _RAND_607 = {1{`RANDOM}};
  pipe_b_47_1 = _RAND_607[19:0];
  _RAND_608 = {1{`RANDOM}};
  pipe_b_48_0 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  pipe_b_48_1 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  pipe_b_49_0 = _RAND_610[19:0];
  _RAND_611 = {1{`RANDOM}};
  pipe_b_49_1 = _RAND_611[19:0];
  _RAND_612 = {1{`RANDOM}};
  pipe_b_50_0 = _RAND_612[19:0];
  _RAND_613 = {1{`RANDOM}};
  pipe_b_50_1 = _RAND_613[19:0];
  _RAND_614 = {1{`RANDOM}};
  pipe_b_51_0 = _RAND_614[19:0];
  _RAND_615 = {1{`RANDOM}};
  pipe_b_51_1 = _RAND_615[19:0];
  _RAND_616 = {1{`RANDOM}};
  pipe_b_52_0 = _RAND_616[19:0];
  _RAND_617 = {1{`RANDOM}};
  pipe_b_52_1 = _RAND_617[19:0];
  _RAND_618 = {1{`RANDOM}};
  pipe_b_53_0 = _RAND_618[19:0];
  _RAND_619 = {1{`RANDOM}};
  pipe_b_53_1 = _RAND_619[19:0];
  _RAND_620 = {1{`RANDOM}};
  pipe_b_54_0 = _RAND_620[19:0];
  _RAND_621 = {1{`RANDOM}};
  pipe_b_54_1 = _RAND_621[19:0];
  _RAND_622 = {1{`RANDOM}};
  pipe_b_55_0 = _RAND_622[19:0];
  _RAND_623 = {1{`RANDOM}};
  pipe_b_55_1 = _RAND_623[19:0];
  _RAND_624 = {1{`RANDOM}};
  pipe_b_56_0 = _RAND_624[19:0];
  _RAND_625 = {1{`RANDOM}};
  pipe_b_56_1 = _RAND_625[19:0];
  _RAND_626 = {1{`RANDOM}};
  pipe_b_57_0 = _RAND_626[19:0];
  _RAND_627 = {1{`RANDOM}};
  pipe_b_57_1 = _RAND_627[19:0];
  _RAND_628 = {1{`RANDOM}};
  pipe_b_58_0 = _RAND_628[19:0];
  _RAND_629 = {1{`RANDOM}};
  pipe_b_58_1 = _RAND_629[19:0];
  _RAND_630 = {1{`RANDOM}};
  pipe_b_59_0 = _RAND_630[19:0];
  _RAND_631 = {1{`RANDOM}};
  pipe_b_59_1 = _RAND_631[19:0];
  _RAND_632 = {1{`RANDOM}};
  pipe_b_60_0 = _RAND_632[19:0];
  _RAND_633 = {1{`RANDOM}};
  pipe_b_60_1 = _RAND_633[19:0];
  _RAND_634 = {1{`RANDOM}};
  pipe_b_61_0 = _RAND_634[19:0];
  _RAND_635 = {1{`RANDOM}};
  pipe_b_61_1 = _RAND_635[19:0];
  _RAND_636 = {1{`RANDOM}};
  pipe_b_62_0 = _RAND_636[19:0];
  _RAND_637 = {1{`RANDOM}};
  pipe_b_62_1 = _RAND_637[19:0];
  _RAND_638 = {1{`RANDOM}};
  pipe_b_63_0 = _RAND_638[19:0];
  _RAND_639 = {1{`RANDOM}};
  pipe_b_63_1 = _RAND_639[19:0];
  _RAND_640 = {1{`RANDOM}};
  pipe_b_64_0 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  pipe_b_64_1 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  pipe_b_65_0 = _RAND_642[19:0];
  _RAND_643 = {1{`RANDOM}};
  pipe_b_65_1 = _RAND_643[19:0];
  _RAND_644 = {1{`RANDOM}};
  pipe_b_66_0 = _RAND_644[19:0];
  _RAND_645 = {1{`RANDOM}};
  pipe_b_66_1 = _RAND_645[19:0];
  _RAND_646 = {1{`RANDOM}};
  pipe_b_67_0 = _RAND_646[19:0];
  _RAND_647 = {1{`RANDOM}};
  pipe_b_67_1 = _RAND_647[19:0];
  _RAND_648 = {1{`RANDOM}};
  pipe_b_68_0 = _RAND_648[19:0];
  _RAND_649 = {1{`RANDOM}};
  pipe_b_68_1 = _RAND_649[19:0];
  _RAND_650 = {1{`RANDOM}};
  pipe_b_69_0 = _RAND_650[19:0];
  _RAND_651 = {1{`RANDOM}};
  pipe_b_69_1 = _RAND_651[19:0];
  _RAND_652 = {1{`RANDOM}};
  pipe_b_70_0 = _RAND_652[19:0];
  _RAND_653 = {1{`RANDOM}};
  pipe_b_70_1 = _RAND_653[19:0];
  _RAND_654 = {1{`RANDOM}};
  pipe_b_71_0 = _RAND_654[19:0];
  _RAND_655 = {1{`RANDOM}};
  pipe_b_71_1 = _RAND_655[19:0];
  _RAND_656 = {1{`RANDOM}};
  pipe_b_72_0 = _RAND_656[19:0];
  _RAND_657 = {1{`RANDOM}};
  pipe_b_72_1 = _RAND_657[19:0];
  _RAND_658 = {1{`RANDOM}};
  pipe_b_73_0 = _RAND_658[19:0];
  _RAND_659 = {1{`RANDOM}};
  pipe_b_73_1 = _RAND_659[19:0];
  _RAND_660 = {1{`RANDOM}};
  pipe_b_74_0 = _RAND_660[19:0];
  _RAND_661 = {1{`RANDOM}};
  pipe_b_74_1 = _RAND_661[19:0];
  _RAND_662 = {1{`RANDOM}};
  pipe_b_75_0 = _RAND_662[19:0];
  _RAND_663 = {1{`RANDOM}};
  pipe_b_75_1 = _RAND_663[19:0];
  _RAND_664 = {1{`RANDOM}};
  pipe_b_76_0 = _RAND_664[19:0];
  _RAND_665 = {1{`RANDOM}};
  pipe_b_76_1 = _RAND_665[19:0];
  _RAND_666 = {1{`RANDOM}};
  pipe_b_77_0 = _RAND_666[19:0];
  _RAND_667 = {1{`RANDOM}};
  pipe_b_77_1 = _RAND_667[19:0];
  _RAND_668 = {1{`RANDOM}};
  pipe_b_78_0 = _RAND_668[19:0];
  _RAND_669 = {1{`RANDOM}};
  pipe_b_78_1 = _RAND_669[19:0];
  _RAND_670 = {1{`RANDOM}};
  pipe_b_79_0 = _RAND_670[19:0];
  _RAND_671 = {1{`RANDOM}};
  pipe_b_79_1 = _RAND_671[19:0];
  _RAND_672 = {1{`RANDOM}};
  pipe_b_80_0 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  pipe_b_80_1 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  pipe_b_81_0 = _RAND_674[19:0];
  _RAND_675 = {1{`RANDOM}};
  pipe_b_81_1 = _RAND_675[19:0];
  _RAND_676 = {1{`RANDOM}};
  pipe_b_82_0 = _RAND_676[19:0];
  _RAND_677 = {1{`RANDOM}};
  pipe_b_82_1 = _RAND_677[19:0];
  _RAND_678 = {1{`RANDOM}};
  pipe_b_83_0 = _RAND_678[19:0];
  _RAND_679 = {1{`RANDOM}};
  pipe_b_83_1 = _RAND_679[19:0];
  _RAND_680 = {1{`RANDOM}};
  pipe_b_84_0 = _RAND_680[19:0];
  _RAND_681 = {1{`RANDOM}};
  pipe_b_84_1 = _RAND_681[19:0];
  _RAND_682 = {1{`RANDOM}};
  pipe_b_85_0 = _RAND_682[19:0];
  _RAND_683 = {1{`RANDOM}};
  pipe_b_85_1 = _RAND_683[19:0];
  _RAND_684 = {1{`RANDOM}};
  pipe_b_86_0 = _RAND_684[19:0];
  _RAND_685 = {1{`RANDOM}};
  pipe_b_86_1 = _RAND_685[19:0];
  _RAND_686 = {1{`RANDOM}};
  pipe_b_87_0 = _RAND_686[19:0];
  _RAND_687 = {1{`RANDOM}};
  pipe_b_87_1 = _RAND_687[19:0];
  _RAND_688 = {1{`RANDOM}};
  pipe_b_88_0 = _RAND_688[19:0];
  _RAND_689 = {1{`RANDOM}};
  pipe_b_88_1 = _RAND_689[19:0];
  _RAND_690 = {1{`RANDOM}};
  pipe_b_89_0 = _RAND_690[19:0];
  _RAND_691 = {1{`RANDOM}};
  pipe_b_89_1 = _RAND_691[19:0];
  _RAND_692 = {1{`RANDOM}};
  pipe_b_90_0 = _RAND_692[19:0];
  _RAND_693 = {1{`RANDOM}};
  pipe_b_90_1 = _RAND_693[19:0];
  _RAND_694 = {1{`RANDOM}};
  pipe_b_91_0 = _RAND_694[19:0];
  _RAND_695 = {1{`RANDOM}};
  pipe_b_91_1 = _RAND_695[19:0];
  _RAND_696 = {1{`RANDOM}};
  pipe_b_92_0 = _RAND_696[19:0];
  _RAND_697 = {1{`RANDOM}};
  pipe_b_92_1 = _RAND_697[19:0];
  _RAND_698 = {1{`RANDOM}};
  pipe_b_93_0 = _RAND_698[19:0];
  _RAND_699 = {1{`RANDOM}};
  pipe_b_93_1 = _RAND_699[19:0];
  _RAND_700 = {1{`RANDOM}};
  pipe_b_94_0 = _RAND_700[19:0];
  _RAND_701 = {1{`RANDOM}};
  pipe_b_94_1 = _RAND_701[19:0];
  _RAND_702 = {1{`RANDOM}};
  pipe_b_95_0 = _RAND_702[19:0];
  _RAND_703 = {1{`RANDOM}};
  pipe_b_95_1 = _RAND_703[19:0];
  _RAND_704 = {1{`RANDOM}};
  pipe_b_96_0 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  pipe_b_96_1 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  pipe_b_97_0 = _RAND_706[19:0];
  _RAND_707 = {1{`RANDOM}};
  pipe_b_97_1 = _RAND_707[19:0];
  _RAND_708 = {1{`RANDOM}};
  pipe_b_98_0 = _RAND_708[19:0];
  _RAND_709 = {1{`RANDOM}};
  pipe_b_98_1 = _RAND_709[19:0];
  _RAND_710 = {1{`RANDOM}};
  pipe_b_99_0 = _RAND_710[19:0];
  _RAND_711 = {1{`RANDOM}};
  pipe_b_99_1 = _RAND_711[19:0];
  _RAND_712 = {1{`RANDOM}};
  pipe_b_100_0 = _RAND_712[19:0];
  _RAND_713 = {1{`RANDOM}};
  pipe_b_100_1 = _RAND_713[19:0];
  _RAND_714 = {1{`RANDOM}};
  pipe_b_101_0 = _RAND_714[19:0];
  _RAND_715 = {1{`RANDOM}};
  pipe_b_101_1 = _RAND_715[19:0];
  _RAND_716 = {1{`RANDOM}};
  pipe_b_102_0 = _RAND_716[19:0];
  _RAND_717 = {1{`RANDOM}};
  pipe_b_102_1 = _RAND_717[19:0];
  _RAND_718 = {1{`RANDOM}};
  pipe_b_103_0 = _RAND_718[19:0];
  _RAND_719 = {1{`RANDOM}};
  pipe_b_103_1 = _RAND_719[19:0];
  _RAND_720 = {1{`RANDOM}};
  pipe_b_104_0 = _RAND_720[19:0];
  _RAND_721 = {1{`RANDOM}};
  pipe_b_104_1 = _RAND_721[19:0];
  _RAND_722 = {1{`RANDOM}};
  pipe_b_105_0 = _RAND_722[19:0];
  _RAND_723 = {1{`RANDOM}};
  pipe_b_105_1 = _RAND_723[19:0];
  _RAND_724 = {1{`RANDOM}};
  pipe_b_106_0 = _RAND_724[19:0];
  _RAND_725 = {1{`RANDOM}};
  pipe_b_106_1 = _RAND_725[19:0];
  _RAND_726 = {1{`RANDOM}};
  pipe_b_107_0 = _RAND_726[19:0];
  _RAND_727 = {1{`RANDOM}};
  pipe_b_107_1 = _RAND_727[19:0];
  _RAND_728 = {1{`RANDOM}};
  pipe_b_108_0 = _RAND_728[19:0];
  _RAND_729 = {1{`RANDOM}};
  pipe_b_108_1 = _RAND_729[19:0];
  _RAND_730 = {1{`RANDOM}};
  pipe_b_109_0 = _RAND_730[19:0];
  _RAND_731 = {1{`RANDOM}};
  pipe_b_109_1 = _RAND_731[19:0];
  _RAND_732 = {1{`RANDOM}};
  pipe_b_110_0 = _RAND_732[19:0];
  _RAND_733 = {1{`RANDOM}};
  pipe_b_110_1 = _RAND_733[19:0];
  _RAND_734 = {1{`RANDOM}};
  pipe_b_111_0 = _RAND_734[19:0];
  _RAND_735 = {1{`RANDOM}};
  pipe_b_111_1 = _RAND_735[19:0];
  _RAND_736 = {1{`RANDOM}};
  pipe_b_112_0 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  pipe_b_112_1 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  pipe_b_113_0 = _RAND_738[19:0];
  _RAND_739 = {1{`RANDOM}};
  pipe_b_113_1 = _RAND_739[19:0];
  _RAND_740 = {1{`RANDOM}};
  pipe_b_114_0 = _RAND_740[19:0];
  _RAND_741 = {1{`RANDOM}};
  pipe_b_114_1 = _RAND_741[19:0];
  _RAND_742 = {1{`RANDOM}};
  pipe_b_115_0 = _RAND_742[19:0];
  _RAND_743 = {1{`RANDOM}};
  pipe_b_115_1 = _RAND_743[19:0];
  _RAND_744 = {1{`RANDOM}};
  pipe_b_116_0 = _RAND_744[19:0];
  _RAND_745 = {1{`RANDOM}};
  pipe_b_116_1 = _RAND_745[19:0];
  _RAND_746 = {1{`RANDOM}};
  pipe_b_117_0 = _RAND_746[19:0];
  _RAND_747 = {1{`RANDOM}};
  pipe_b_117_1 = _RAND_747[19:0];
  _RAND_748 = {1{`RANDOM}};
  pipe_b_118_0 = _RAND_748[19:0];
  _RAND_749 = {1{`RANDOM}};
  pipe_b_118_1 = _RAND_749[19:0];
  _RAND_750 = {1{`RANDOM}};
  pipe_b_119_0 = _RAND_750[19:0];
  _RAND_751 = {1{`RANDOM}};
  pipe_b_119_1 = _RAND_751[19:0];
  _RAND_752 = {1{`RANDOM}};
  pipe_b_120_0 = _RAND_752[19:0];
  _RAND_753 = {1{`RANDOM}};
  pipe_b_120_1 = _RAND_753[19:0];
  _RAND_754 = {1{`RANDOM}};
  pipe_b_121_0 = _RAND_754[19:0];
  _RAND_755 = {1{`RANDOM}};
  pipe_b_121_1 = _RAND_755[19:0];
  _RAND_756 = {1{`RANDOM}};
  pipe_b_122_0 = _RAND_756[19:0];
  _RAND_757 = {1{`RANDOM}};
  pipe_b_122_1 = _RAND_757[19:0];
  _RAND_758 = {1{`RANDOM}};
  pipe_b_123_0 = _RAND_758[19:0];
  _RAND_759 = {1{`RANDOM}};
  pipe_b_123_1 = _RAND_759[19:0];
  _RAND_760 = {1{`RANDOM}};
  pipe_b_124_0 = _RAND_760[19:0];
  _RAND_761 = {1{`RANDOM}};
  pipe_b_124_1 = _RAND_761[19:0];
  _RAND_762 = {1{`RANDOM}};
  pipe_b_125_0 = _RAND_762[19:0];
  _RAND_763 = {1{`RANDOM}};
  pipe_b_125_1 = _RAND_763[19:0];
  _RAND_764 = {1{`RANDOM}};
  pipe_b_126_0 = _RAND_764[19:0];
  _RAND_765 = {1{`RANDOM}};
  pipe_b_126_1 = _RAND_765[19:0];
  _RAND_766 = {1{`RANDOM}};
  pipe_b_127_0 = _RAND_766[19:0];
  _RAND_767 = {1{`RANDOM}};
  pipe_b_127_1 = _RAND_767[19:0];
  _RAND_768 = {1{`RANDOM}};
  pipe_b_128_0 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  pipe_b_128_1 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  pipe_b_129_0 = _RAND_770[19:0];
  _RAND_771 = {1{`RANDOM}};
  pipe_b_129_1 = _RAND_771[19:0];
  _RAND_772 = {1{`RANDOM}};
  pipe_b_130_0 = _RAND_772[19:0];
  _RAND_773 = {1{`RANDOM}};
  pipe_b_130_1 = _RAND_773[19:0];
  _RAND_774 = {1{`RANDOM}};
  pipe_b_131_0 = _RAND_774[19:0];
  _RAND_775 = {1{`RANDOM}};
  pipe_b_131_1 = _RAND_775[19:0];
  _RAND_776 = {1{`RANDOM}};
  pipe_b_132_0 = _RAND_776[19:0];
  _RAND_777 = {1{`RANDOM}};
  pipe_b_132_1 = _RAND_777[19:0];
  _RAND_778 = {1{`RANDOM}};
  pipe_b_133_0 = _RAND_778[19:0];
  _RAND_779 = {1{`RANDOM}};
  pipe_b_133_1 = _RAND_779[19:0];
  _RAND_780 = {1{`RANDOM}};
  pipe_b_134_0 = _RAND_780[19:0];
  _RAND_781 = {1{`RANDOM}};
  pipe_b_134_1 = _RAND_781[19:0];
  _RAND_782 = {1{`RANDOM}};
  pipe_b_135_0 = _RAND_782[19:0];
  _RAND_783 = {1{`RANDOM}};
  pipe_b_135_1 = _RAND_783[19:0];
  _RAND_784 = {1{`RANDOM}};
  pipe_b_136_0 = _RAND_784[19:0];
  _RAND_785 = {1{`RANDOM}};
  pipe_b_136_1 = _RAND_785[19:0];
  _RAND_786 = {1{`RANDOM}};
  pipe_b_137_0 = _RAND_786[19:0];
  _RAND_787 = {1{`RANDOM}};
  pipe_b_137_1 = _RAND_787[19:0];
  _RAND_788 = {1{`RANDOM}};
  pipe_b_138_0 = _RAND_788[19:0];
  _RAND_789 = {1{`RANDOM}};
  pipe_b_138_1 = _RAND_789[19:0];
  _RAND_790 = {1{`RANDOM}};
  pipe_b_139_0 = _RAND_790[19:0];
  _RAND_791 = {1{`RANDOM}};
  pipe_b_139_1 = _RAND_791[19:0];
  _RAND_792 = {1{`RANDOM}};
  pipe_b_140_0 = _RAND_792[19:0];
  _RAND_793 = {1{`RANDOM}};
  pipe_b_140_1 = _RAND_793[19:0];
  _RAND_794 = {1{`RANDOM}};
  pipe_b_141_0 = _RAND_794[19:0];
  _RAND_795 = {1{`RANDOM}};
  pipe_b_141_1 = _RAND_795[19:0];
  _RAND_796 = {1{`RANDOM}};
  pipe_b_142_0 = _RAND_796[19:0];
  _RAND_797 = {1{`RANDOM}};
  pipe_b_142_1 = _RAND_797[19:0];
  _RAND_798 = {1{`RANDOM}};
  pipe_b_143_0 = _RAND_798[19:0];
  _RAND_799 = {1{`RANDOM}};
  pipe_b_143_1 = _RAND_799[19:0];
  _RAND_800 = {1{`RANDOM}};
  pipe_b_144_0 = _RAND_800[7:0];
  _RAND_801 = {1{`RANDOM}};
  pipe_b_144_1 = _RAND_801[7:0];
  _RAND_802 = {1{`RANDOM}};
  pipe_b_145_0 = _RAND_802[19:0];
  _RAND_803 = {1{`RANDOM}};
  pipe_b_145_1 = _RAND_803[19:0];
  _RAND_804 = {1{`RANDOM}};
  pipe_b_146_0 = _RAND_804[19:0];
  _RAND_805 = {1{`RANDOM}};
  pipe_b_146_1 = _RAND_805[19:0];
  _RAND_806 = {1{`RANDOM}};
  pipe_b_147_0 = _RAND_806[19:0];
  _RAND_807 = {1{`RANDOM}};
  pipe_b_147_1 = _RAND_807[19:0];
  _RAND_808 = {1{`RANDOM}};
  pipe_b_148_0 = _RAND_808[19:0];
  _RAND_809 = {1{`RANDOM}};
  pipe_b_148_1 = _RAND_809[19:0];
  _RAND_810 = {1{`RANDOM}};
  pipe_b_149_0 = _RAND_810[19:0];
  _RAND_811 = {1{`RANDOM}};
  pipe_b_149_1 = _RAND_811[19:0];
  _RAND_812 = {1{`RANDOM}};
  pipe_b_150_0 = _RAND_812[19:0];
  _RAND_813 = {1{`RANDOM}};
  pipe_b_150_1 = _RAND_813[19:0];
  _RAND_814 = {1{`RANDOM}};
  pipe_b_151_0 = _RAND_814[19:0];
  _RAND_815 = {1{`RANDOM}};
  pipe_b_151_1 = _RAND_815[19:0];
  _RAND_816 = {1{`RANDOM}};
  pipe_b_152_0 = _RAND_816[19:0];
  _RAND_817 = {1{`RANDOM}};
  pipe_b_152_1 = _RAND_817[19:0];
  _RAND_818 = {1{`RANDOM}};
  pipe_b_153_0 = _RAND_818[19:0];
  _RAND_819 = {1{`RANDOM}};
  pipe_b_153_1 = _RAND_819[19:0];
  _RAND_820 = {1{`RANDOM}};
  pipe_b_154_0 = _RAND_820[19:0];
  _RAND_821 = {1{`RANDOM}};
  pipe_b_154_1 = _RAND_821[19:0];
  _RAND_822 = {1{`RANDOM}};
  pipe_b_155_0 = _RAND_822[19:0];
  _RAND_823 = {1{`RANDOM}};
  pipe_b_155_1 = _RAND_823[19:0];
  _RAND_824 = {1{`RANDOM}};
  pipe_b_156_0 = _RAND_824[19:0];
  _RAND_825 = {1{`RANDOM}};
  pipe_b_156_1 = _RAND_825[19:0];
  _RAND_826 = {1{`RANDOM}};
  pipe_b_157_0 = _RAND_826[19:0];
  _RAND_827 = {1{`RANDOM}};
  pipe_b_157_1 = _RAND_827[19:0];
  _RAND_828 = {1{`RANDOM}};
  pipe_b_158_0 = _RAND_828[19:0];
  _RAND_829 = {1{`RANDOM}};
  pipe_b_158_1 = _RAND_829[19:0];
  _RAND_830 = {1{`RANDOM}};
  pipe_b_159_0 = _RAND_830[19:0];
  _RAND_831 = {1{`RANDOM}};
  pipe_b_159_1 = _RAND_831[19:0];
  _RAND_832 = {1{`RANDOM}};
  pipe_b_160_0 = _RAND_832[7:0];
  _RAND_833 = {1{`RANDOM}};
  pipe_b_160_1 = _RAND_833[7:0];
  _RAND_834 = {1{`RANDOM}};
  pipe_b_161_0 = _RAND_834[19:0];
  _RAND_835 = {1{`RANDOM}};
  pipe_b_161_1 = _RAND_835[19:0];
  _RAND_836 = {1{`RANDOM}};
  pipe_b_162_0 = _RAND_836[19:0];
  _RAND_837 = {1{`RANDOM}};
  pipe_b_162_1 = _RAND_837[19:0];
  _RAND_838 = {1{`RANDOM}};
  pipe_b_163_0 = _RAND_838[19:0];
  _RAND_839 = {1{`RANDOM}};
  pipe_b_163_1 = _RAND_839[19:0];
  _RAND_840 = {1{`RANDOM}};
  pipe_b_164_0 = _RAND_840[19:0];
  _RAND_841 = {1{`RANDOM}};
  pipe_b_164_1 = _RAND_841[19:0];
  _RAND_842 = {1{`RANDOM}};
  pipe_b_165_0 = _RAND_842[19:0];
  _RAND_843 = {1{`RANDOM}};
  pipe_b_165_1 = _RAND_843[19:0];
  _RAND_844 = {1{`RANDOM}};
  pipe_b_166_0 = _RAND_844[19:0];
  _RAND_845 = {1{`RANDOM}};
  pipe_b_166_1 = _RAND_845[19:0];
  _RAND_846 = {1{`RANDOM}};
  pipe_b_167_0 = _RAND_846[19:0];
  _RAND_847 = {1{`RANDOM}};
  pipe_b_167_1 = _RAND_847[19:0];
  _RAND_848 = {1{`RANDOM}};
  pipe_b_168_0 = _RAND_848[19:0];
  _RAND_849 = {1{`RANDOM}};
  pipe_b_168_1 = _RAND_849[19:0];
  _RAND_850 = {1{`RANDOM}};
  pipe_b_169_0 = _RAND_850[19:0];
  _RAND_851 = {1{`RANDOM}};
  pipe_b_169_1 = _RAND_851[19:0];
  _RAND_852 = {1{`RANDOM}};
  pipe_b_170_0 = _RAND_852[19:0];
  _RAND_853 = {1{`RANDOM}};
  pipe_b_170_1 = _RAND_853[19:0];
  _RAND_854 = {1{`RANDOM}};
  pipe_b_171_0 = _RAND_854[19:0];
  _RAND_855 = {1{`RANDOM}};
  pipe_b_171_1 = _RAND_855[19:0];
  _RAND_856 = {1{`RANDOM}};
  pipe_b_172_0 = _RAND_856[19:0];
  _RAND_857 = {1{`RANDOM}};
  pipe_b_172_1 = _RAND_857[19:0];
  _RAND_858 = {1{`RANDOM}};
  pipe_b_173_0 = _RAND_858[19:0];
  _RAND_859 = {1{`RANDOM}};
  pipe_b_173_1 = _RAND_859[19:0];
  _RAND_860 = {1{`RANDOM}};
  pipe_b_174_0 = _RAND_860[19:0];
  _RAND_861 = {1{`RANDOM}};
  pipe_b_174_1 = _RAND_861[19:0];
  _RAND_862 = {1{`RANDOM}};
  pipe_b_175_0 = _RAND_862[19:0];
  _RAND_863 = {1{`RANDOM}};
  pipe_b_175_1 = _RAND_863[19:0];
  _RAND_864 = {1{`RANDOM}};
  pipe_b_176_0 = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  pipe_b_176_1 = _RAND_865[7:0];
  _RAND_866 = {1{`RANDOM}};
  pipe_b_177_0 = _RAND_866[19:0];
  _RAND_867 = {1{`RANDOM}};
  pipe_b_177_1 = _RAND_867[19:0];
  _RAND_868 = {1{`RANDOM}};
  pipe_b_178_0 = _RAND_868[19:0];
  _RAND_869 = {1{`RANDOM}};
  pipe_b_178_1 = _RAND_869[19:0];
  _RAND_870 = {1{`RANDOM}};
  pipe_b_179_0 = _RAND_870[19:0];
  _RAND_871 = {1{`RANDOM}};
  pipe_b_179_1 = _RAND_871[19:0];
  _RAND_872 = {1{`RANDOM}};
  pipe_b_180_0 = _RAND_872[19:0];
  _RAND_873 = {1{`RANDOM}};
  pipe_b_180_1 = _RAND_873[19:0];
  _RAND_874 = {1{`RANDOM}};
  pipe_b_181_0 = _RAND_874[19:0];
  _RAND_875 = {1{`RANDOM}};
  pipe_b_181_1 = _RAND_875[19:0];
  _RAND_876 = {1{`RANDOM}};
  pipe_b_182_0 = _RAND_876[19:0];
  _RAND_877 = {1{`RANDOM}};
  pipe_b_182_1 = _RAND_877[19:0];
  _RAND_878 = {1{`RANDOM}};
  pipe_b_183_0 = _RAND_878[19:0];
  _RAND_879 = {1{`RANDOM}};
  pipe_b_183_1 = _RAND_879[19:0];
  _RAND_880 = {1{`RANDOM}};
  pipe_b_184_0 = _RAND_880[19:0];
  _RAND_881 = {1{`RANDOM}};
  pipe_b_184_1 = _RAND_881[19:0];
  _RAND_882 = {1{`RANDOM}};
  pipe_b_185_0 = _RAND_882[19:0];
  _RAND_883 = {1{`RANDOM}};
  pipe_b_185_1 = _RAND_883[19:0];
  _RAND_884 = {1{`RANDOM}};
  pipe_b_186_0 = _RAND_884[19:0];
  _RAND_885 = {1{`RANDOM}};
  pipe_b_186_1 = _RAND_885[19:0];
  _RAND_886 = {1{`RANDOM}};
  pipe_b_187_0 = _RAND_886[19:0];
  _RAND_887 = {1{`RANDOM}};
  pipe_b_187_1 = _RAND_887[19:0];
  _RAND_888 = {1{`RANDOM}};
  pipe_b_188_0 = _RAND_888[19:0];
  _RAND_889 = {1{`RANDOM}};
  pipe_b_188_1 = _RAND_889[19:0];
  _RAND_890 = {1{`RANDOM}};
  pipe_b_189_0 = _RAND_890[19:0];
  _RAND_891 = {1{`RANDOM}};
  pipe_b_189_1 = _RAND_891[19:0];
  _RAND_892 = {1{`RANDOM}};
  pipe_b_190_0 = _RAND_892[19:0];
  _RAND_893 = {1{`RANDOM}};
  pipe_b_190_1 = _RAND_893[19:0];
  _RAND_894 = {1{`RANDOM}};
  pipe_b_191_0 = _RAND_894[19:0];
  _RAND_895 = {1{`RANDOM}};
  pipe_b_191_1 = _RAND_895[19:0];
  _RAND_896 = {1{`RANDOM}};
  pipe_b_192_0 = _RAND_896[7:0];
  _RAND_897 = {1{`RANDOM}};
  pipe_b_192_1 = _RAND_897[7:0];
  _RAND_898 = {1{`RANDOM}};
  pipe_b_193_0 = _RAND_898[19:0];
  _RAND_899 = {1{`RANDOM}};
  pipe_b_193_1 = _RAND_899[19:0];
  _RAND_900 = {1{`RANDOM}};
  pipe_b_194_0 = _RAND_900[19:0];
  _RAND_901 = {1{`RANDOM}};
  pipe_b_194_1 = _RAND_901[19:0];
  _RAND_902 = {1{`RANDOM}};
  pipe_b_195_0 = _RAND_902[19:0];
  _RAND_903 = {1{`RANDOM}};
  pipe_b_195_1 = _RAND_903[19:0];
  _RAND_904 = {1{`RANDOM}};
  pipe_b_196_0 = _RAND_904[19:0];
  _RAND_905 = {1{`RANDOM}};
  pipe_b_196_1 = _RAND_905[19:0];
  _RAND_906 = {1{`RANDOM}};
  pipe_b_197_0 = _RAND_906[19:0];
  _RAND_907 = {1{`RANDOM}};
  pipe_b_197_1 = _RAND_907[19:0];
  _RAND_908 = {1{`RANDOM}};
  pipe_b_198_0 = _RAND_908[19:0];
  _RAND_909 = {1{`RANDOM}};
  pipe_b_198_1 = _RAND_909[19:0];
  _RAND_910 = {1{`RANDOM}};
  pipe_b_199_0 = _RAND_910[19:0];
  _RAND_911 = {1{`RANDOM}};
  pipe_b_199_1 = _RAND_911[19:0];
  _RAND_912 = {1{`RANDOM}};
  pipe_b_200_0 = _RAND_912[19:0];
  _RAND_913 = {1{`RANDOM}};
  pipe_b_200_1 = _RAND_913[19:0];
  _RAND_914 = {1{`RANDOM}};
  pipe_b_201_0 = _RAND_914[19:0];
  _RAND_915 = {1{`RANDOM}};
  pipe_b_201_1 = _RAND_915[19:0];
  _RAND_916 = {1{`RANDOM}};
  pipe_b_202_0 = _RAND_916[19:0];
  _RAND_917 = {1{`RANDOM}};
  pipe_b_202_1 = _RAND_917[19:0];
  _RAND_918 = {1{`RANDOM}};
  pipe_b_203_0 = _RAND_918[19:0];
  _RAND_919 = {1{`RANDOM}};
  pipe_b_203_1 = _RAND_919[19:0];
  _RAND_920 = {1{`RANDOM}};
  pipe_b_204_0 = _RAND_920[19:0];
  _RAND_921 = {1{`RANDOM}};
  pipe_b_204_1 = _RAND_921[19:0];
  _RAND_922 = {1{`RANDOM}};
  pipe_b_205_0 = _RAND_922[19:0];
  _RAND_923 = {1{`RANDOM}};
  pipe_b_205_1 = _RAND_923[19:0];
  _RAND_924 = {1{`RANDOM}};
  pipe_b_206_0 = _RAND_924[19:0];
  _RAND_925 = {1{`RANDOM}};
  pipe_b_206_1 = _RAND_925[19:0];
  _RAND_926 = {1{`RANDOM}};
  pipe_b_207_0 = _RAND_926[19:0];
  _RAND_927 = {1{`RANDOM}};
  pipe_b_207_1 = _RAND_927[19:0];
  _RAND_928 = {1{`RANDOM}};
  pipe_b_208_0 = _RAND_928[7:0];
  _RAND_929 = {1{`RANDOM}};
  pipe_b_208_1 = _RAND_929[7:0];
  _RAND_930 = {1{`RANDOM}};
  pipe_b_209_0 = _RAND_930[19:0];
  _RAND_931 = {1{`RANDOM}};
  pipe_b_209_1 = _RAND_931[19:0];
  _RAND_932 = {1{`RANDOM}};
  pipe_b_210_0 = _RAND_932[19:0];
  _RAND_933 = {1{`RANDOM}};
  pipe_b_210_1 = _RAND_933[19:0];
  _RAND_934 = {1{`RANDOM}};
  pipe_b_211_0 = _RAND_934[19:0];
  _RAND_935 = {1{`RANDOM}};
  pipe_b_211_1 = _RAND_935[19:0];
  _RAND_936 = {1{`RANDOM}};
  pipe_b_212_0 = _RAND_936[19:0];
  _RAND_937 = {1{`RANDOM}};
  pipe_b_212_1 = _RAND_937[19:0];
  _RAND_938 = {1{`RANDOM}};
  pipe_b_213_0 = _RAND_938[19:0];
  _RAND_939 = {1{`RANDOM}};
  pipe_b_213_1 = _RAND_939[19:0];
  _RAND_940 = {1{`RANDOM}};
  pipe_b_214_0 = _RAND_940[19:0];
  _RAND_941 = {1{`RANDOM}};
  pipe_b_214_1 = _RAND_941[19:0];
  _RAND_942 = {1{`RANDOM}};
  pipe_b_215_0 = _RAND_942[19:0];
  _RAND_943 = {1{`RANDOM}};
  pipe_b_215_1 = _RAND_943[19:0];
  _RAND_944 = {1{`RANDOM}};
  pipe_b_216_0 = _RAND_944[19:0];
  _RAND_945 = {1{`RANDOM}};
  pipe_b_216_1 = _RAND_945[19:0];
  _RAND_946 = {1{`RANDOM}};
  pipe_b_217_0 = _RAND_946[19:0];
  _RAND_947 = {1{`RANDOM}};
  pipe_b_217_1 = _RAND_947[19:0];
  _RAND_948 = {1{`RANDOM}};
  pipe_b_218_0 = _RAND_948[19:0];
  _RAND_949 = {1{`RANDOM}};
  pipe_b_218_1 = _RAND_949[19:0];
  _RAND_950 = {1{`RANDOM}};
  pipe_b_219_0 = _RAND_950[19:0];
  _RAND_951 = {1{`RANDOM}};
  pipe_b_219_1 = _RAND_951[19:0];
  _RAND_952 = {1{`RANDOM}};
  pipe_b_220_0 = _RAND_952[19:0];
  _RAND_953 = {1{`RANDOM}};
  pipe_b_220_1 = _RAND_953[19:0];
  _RAND_954 = {1{`RANDOM}};
  pipe_b_221_0 = _RAND_954[19:0];
  _RAND_955 = {1{`RANDOM}};
  pipe_b_221_1 = _RAND_955[19:0];
  _RAND_956 = {1{`RANDOM}};
  pipe_b_222_0 = _RAND_956[19:0];
  _RAND_957 = {1{`RANDOM}};
  pipe_b_222_1 = _RAND_957[19:0];
  _RAND_958 = {1{`RANDOM}};
  pipe_b_223_0 = _RAND_958[19:0];
  _RAND_959 = {1{`RANDOM}};
  pipe_b_223_1 = _RAND_959[19:0];
  _RAND_960 = {1{`RANDOM}};
  pipe_b_224_0 = _RAND_960[7:0];
  _RAND_961 = {1{`RANDOM}};
  pipe_b_224_1 = _RAND_961[7:0];
  _RAND_962 = {1{`RANDOM}};
  pipe_b_225_0 = _RAND_962[19:0];
  _RAND_963 = {1{`RANDOM}};
  pipe_b_225_1 = _RAND_963[19:0];
  _RAND_964 = {1{`RANDOM}};
  pipe_b_226_0 = _RAND_964[19:0];
  _RAND_965 = {1{`RANDOM}};
  pipe_b_226_1 = _RAND_965[19:0];
  _RAND_966 = {1{`RANDOM}};
  pipe_b_227_0 = _RAND_966[19:0];
  _RAND_967 = {1{`RANDOM}};
  pipe_b_227_1 = _RAND_967[19:0];
  _RAND_968 = {1{`RANDOM}};
  pipe_b_228_0 = _RAND_968[19:0];
  _RAND_969 = {1{`RANDOM}};
  pipe_b_228_1 = _RAND_969[19:0];
  _RAND_970 = {1{`RANDOM}};
  pipe_b_229_0 = _RAND_970[19:0];
  _RAND_971 = {1{`RANDOM}};
  pipe_b_229_1 = _RAND_971[19:0];
  _RAND_972 = {1{`RANDOM}};
  pipe_b_230_0 = _RAND_972[19:0];
  _RAND_973 = {1{`RANDOM}};
  pipe_b_230_1 = _RAND_973[19:0];
  _RAND_974 = {1{`RANDOM}};
  pipe_b_231_0 = _RAND_974[19:0];
  _RAND_975 = {1{`RANDOM}};
  pipe_b_231_1 = _RAND_975[19:0];
  _RAND_976 = {1{`RANDOM}};
  pipe_b_232_0 = _RAND_976[19:0];
  _RAND_977 = {1{`RANDOM}};
  pipe_b_232_1 = _RAND_977[19:0];
  _RAND_978 = {1{`RANDOM}};
  pipe_b_233_0 = _RAND_978[19:0];
  _RAND_979 = {1{`RANDOM}};
  pipe_b_233_1 = _RAND_979[19:0];
  _RAND_980 = {1{`RANDOM}};
  pipe_b_234_0 = _RAND_980[19:0];
  _RAND_981 = {1{`RANDOM}};
  pipe_b_234_1 = _RAND_981[19:0];
  _RAND_982 = {1{`RANDOM}};
  pipe_b_235_0 = _RAND_982[19:0];
  _RAND_983 = {1{`RANDOM}};
  pipe_b_235_1 = _RAND_983[19:0];
  _RAND_984 = {1{`RANDOM}};
  pipe_b_236_0 = _RAND_984[19:0];
  _RAND_985 = {1{`RANDOM}};
  pipe_b_236_1 = _RAND_985[19:0];
  _RAND_986 = {1{`RANDOM}};
  pipe_b_237_0 = _RAND_986[19:0];
  _RAND_987 = {1{`RANDOM}};
  pipe_b_237_1 = _RAND_987[19:0];
  _RAND_988 = {1{`RANDOM}};
  pipe_b_238_0 = _RAND_988[19:0];
  _RAND_989 = {1{`RANDOM}};
  pipe_b_238_1 = _RAND_989[19:0];
  _RAND_990 = {1{`RANDOM}};
  pipe_b_239_0 = _RAND_990[19:0];
  _RAND_991 = {1{`RANDOM}};
  pipe_b_239_1 = _RAND_991[19:0];
  _RAND_992 = {1{`RANDOM}};
  pipe_b_240_0 = _RAND_992[7:0];
  _RAND_993 = {1{`RANDOM}};
  pipe_b_240_1 = _RAND_993[7:0];
  _RAND_994 = {1{`RANDOM}};
  pipe_b_241_0 = _RAND_994[19:0];
  _RAND_995 = {1{`RANDOM}};
  pipe_b_241_1 = _RAND_995[19:0];
  _RAND_996 = {1{`RANDOM}};
  pipe_b_242_0 = _RAND_996[19:0];
  _RAND_997 = {1{`RANDOM}};
  pipe_b_242_1 = _RAND_997[19:0];
  _RAND_998 = {1{`RANDOM}};
  pipe_b_243_0 = _RAND_998[19:0];
  _RAND_999 = {1{`RANDOM}};
  pipe_b_243_1 = _RAND_999[19:0];
  _RAND_1000 = {1{`RANDOM}};
  pipe_b_244_0 = _RAND_1000[19:0];
  _RAND_1001 = {1{`RANDOM}};
  pipe_b_244_1 = _RAND_1001[19:0];
  _RAND_1002 = {1{`RANDOM}};
  pipe_b_245_0 = _RAND_1002[19:0];
  _RAND_1003 = {1{`RANDOM}};
  pipe_b_245_1 = _RAND_1003[19:0];
  _RAND_1004 = {1{`RANDOM}};
  pipe_b_246_0 = _RAND_1004[19:0];
  _RAND_1005 = {1{`RANDOM}};
  pipe_b_246_1 = _RAND_1005[19:0];
  _RAND_1006 = {1{`RANDOM}};
  pipe_b_247_0 = _RAND_1006[19:0];
  _RAND_1007 = {1{`RANDOM}};
  pipe_b_247_1 = _RAND_1007[19:0];
  _RAND_1008 = {1{`RANDOM}};
  pipe_b_248_0 = _RAND_1008[19:0];
  _RAND_1009 = {1{`RANDOM}};
  pipe_b_248_1 = _RAND_1009[19:0];
  _RAND_1010 = {1{`RANDOM}};
  pipe_b_249_0 = _RAND_1010[19:0];
  _RAND_1011 = {1{`RANDOM}};
  pipe_b_249_1 = _RAND_1011[19:0];
  _RAND_1012 = {1{`RANDOM}};
  pipe_b_250_0 = _RAND_1012[19:0];
  _RAND_1013 = {1{`RANDOM}};
  pipe_b_250_1 = _RAND_1013[19:0];
  _RAND_1014 = {1{`RANDOM}};
  pipe_b_251_0 = _RAND_1014[19:0];
  _RAND_1015 = {1{`RANDOM}};
  pipe_b_251_1 = _RAND_1015[19:0];
  _RAND_1016 = {1{`RANDOM}};
  pipe_b_252_0 = _RAND_1016[19:0];
  _RAND_1017 = {1{`RANDOM}};
  pipe_b_252_1 = _RAND_1017[19:0];
  _RAND_1018 = {1{`RANDOM}};
  pipe_b_253_0 = _RAND_1018[19:0];
  _RAND_1019 = {1{`RANDOM}};
  pipe_b_253_1 = _RAND_1019[19:0];
  _RAND_1020 = {1{`RANDOM}};
  pipe_b_254_0 = _RAND_1020[19:0];
  _RAND_1021 = {1{`RANDOM}};
  pipe_b_254_1 = _RAND_1021[19:0];
  _RAND_1022 = {1{`RANDOM}};
  pipe_b_255_0 = _RAND_1022[19:0];
  _RAND_1023 = {1{`RANDOM}};
  pipe_b_255_1 = _RAND_1023[19:0];
  _RAND_1024 = {1{`RANDOM}};
  pipe_b_256_0 = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  pipe_b_256_1 = _RAND_1025[7:0];
  _RAND_1026 = {1{`RANDOM}};
  pipe_b_257_0 = _RAND_1026[19:0];
  _RAND_1027 = {1{`RANDOM}};
  pipe_b_257_1 = _RAND_1027[19:0];
  _RAND_1028 = {1{`RANDOM}};
  pipe_b_258_0 = _RAND_1028[19:0];
  _RAND_1029 = {1{`RANDOM}};
  pipe_b_258_1 = _RAND_1029[19:0];
  _RAND_1030 = {1{`RANDOM}};
  pipe_b_259_0 = _RAND_1030[19:0];
  _RAND_1031 = {1{`RANDOM}};
  pipe_b_259_1 = _RAND_1031[19:0];
  _RAND_1032 = {1{`RANDOM}};
  pipe_b_260_0 = _RAND_1032[19:0];
  _RAND_1033 = {1{`RANDOM}};
  pipe_b_260_1 = _RAND_1033[19:0];
  _RAND_1034 = {1{`RANDOM}};
  pipe_b_261_0 = _RAND_1034[19:0];
  _RAND_1035 = {1{`RANDOM}};
  pipe_b_261_1 = _RAND_1035[19:0];
  _RAND_1036 = {1{`RANDOM}};
  pipe_b_262_0 = _RAND_1036[19:0];
  _RAND_1037 = {1{`RANDOM}};
  pipe_b_262_1 = _RAND_1037[19:0];
  _RAND_1038 = {1{`RANDOM}};
  pipe_b_263_0 = _RAND_1038[19:0];
  _RAND_1039 = {1{`RANDOM}};
  pipe_b_263_1 = _RAND_1039[19:0];
  _RAND_1040 = {1{`RANDOM}};
  pipe_b_264_0 = _RAND_1040[19:0];
  _RAND_1041 = {1{`RANDOM}};
  pipe_b_264_1 = _RAND_1041[19:0];
  _RAND_1042 = {1{`RANDOM}};
  pipe_b_265_0 = _RAND_1042[19:0];
  _RAND_1043 = {1{`RANDOM}};
  pipe_b_265_1 = _RAND_1043[19:0];
  _RAND_1044 = {1{`RANDOM}};
  pipe_b_266_0 = _RAND_1044[19:0];
  _RAND_1045 = {1{`RANDOM}};
  pipe_b_266_1 = _RAND_1045[19:0];
  _RAND_1046 = {1{`RANDOM}};
  pipe_b_267_0 = _RAND_1046[19:0];
  _RAND_1047 = {1{`RANDOM}};
  pipe_b_267_1 = _RAND_1047[19:0];
  _RAND_1048 = {1{`RANDOM}};
  pipe_b_268_0 = _RAND_1048[19:0];
  _RAND_1049 = {1{`RANDOM}};
  pipe_b_268_1 = _RAND_1049[19:0];
  _RAND_1050 = {1{`RANDOM}};
  pipe_b_269_0 = _RAND_1050[19:0];
  _RAND_1051 = {1{`RANDOM}};
  pipe_b_269_1 = _RAND_1051[19:0];
  _RAND_1052 = {1{`RANDOM}};
  pipe_b_270_0 = _RAND_1052[19:0];
  _RAND_1053 = {1{`RANDOM}};
  pipe_b_270_1 = _RAND_1053[19:0];
  _RAND_1054 = {1{`RANDOM}};
  pipe_b_271_0 = _RAND_1054[19:0];
  _RAND_1055 = {1{`RANDOM}};
  pipe_b_271_1 = _RAND_1055[19:0];
  _RAND_1056 = {1{`RANDOM}};
  pipe_b_272_0 = _RAND_1056[7:0];
  _RAND_1057 = {1{`RANDOM}};
  pipe_b_272_1 = _RAND_1057[7:0];
  _RAND_1058 = {1{`RANDOM}};
  pipe_b_273_0 = _RAND_1058[19:0];
  _RAND_1059 = {1{`RANDOM}};
  pipe_b_273_1 = _RAND_1059[19:0];
  _RAND_1060 = {1{`RANDOM}};
  pipe_b_274_0 = _RAND_1060[19:0];
  _RAND_1061 = {1{`RANDOM}};
  pipe_b_274_1 = _RAND_1061[19:0];
  _RAND_1062 = {1{`RANDOM}};
  pipe_b_275_0 = _RAND_1062[19:0];
  _RAND_1063 = {1{`RANDOM}};
  pipe_b_275_1 = _RAND_1063[19:0];
  _RAND_1064 = {1{`RANDOM}};
  pipe_b_276_0 = _RAND_1064[19:0];
  _RAND_1065 = {1{`RANDOM}};
  pipe_b_276_1 = _RAND_1065[19:0];
  _RAND_1066 = {1{`RANDOM}};
  pipe_b_277_0 = _RAND_1066[19:0];
  _RAND_1067 = {1{`RANDOM}};
  pipe_b_277_1 = _RAND_1067[19:0];
  _RAND_1068 = {1{`RANDOM}};
  pipe_b_278_0 = _RAND_1068[19:0];
  _RAND_1069 = {1{`RANDOM}};
  pipe_b_278_1 = _RAND_1069[19:0];
  _RAND_1070 = {1{`RANDOM}};
  pipe_b_279_0 = _RAND_1070[19:0];
  _RAND_1071 = {1{`RANDOM}};
  pipe_b_279_1 = _RAND_1071[19:0];
  _RAND_1072 = {1{`RANDOM}};
  pipe_b_280_0 = _RAND_1072[19:0];
  _RAND_1073 = {1{`RANDOM}};
  pipe_b_280_1 = _RAND_1073[19:0];
  _RAND_1074 = {1{`RANDOM}};
  pipe_b_281_0 = _RAND_1074[19:0];
  _RAND_1075 = {1{`RANDOM}};
  pipe_b_281_1 = _RAND_1075[19:0];
  _RAND_1076 = {1{`RANDOM}};
  pipe_b_282_0 = _RAND_1076[19:0];
  _RAND_1077 = {1{`RANDOM}};
  pipe_b_282_1 = _RAND_1077[19:0];
  _RAND_1078 = {1{`RANDOM}};
  pipe_b_283_0 = _RAND_1078[19:0];
  _RAND_1079 = {1{`RANDOM}};
  pipe_b_283_1 = _RAND_1079[19:0];
  _RAND_1080 = {1{`RANDOM}};
  pipe_b_284_0 = _RAND_1080[19:0];
  _RAND_1081 = {1{`RANDOM}};
  pipe_b_284_1 = _RAND_1081[19:0];
  _RAND_1082 = {1{`RANDOM}};
  pipe_b_285_0 = _RAND_1082[19:0];
  _RAND_1083 = {1{`RANDOM}};
  pipe_b_285_1 = _RAND_1083[19:0];
  _RAND_1084 = {1{`RANDOM}};
  pipe_b_286_0 = _RAND_1084[19:0];
  _RAND_1085 = {1{`RANDOM}};
  pipe_b_286_1 = _RAND_1085[19:0];
  _RAND_1086 = {1{`RANDOM}};
  pipe_b_287_0 = _RAND_1086[19:0];
  _RAND_1087 = {1{`RANDOM}};
  pipe_b_287_1 = _RAND_1087[19:0];
  _RAND_1088 = {1{`RANDOM}};
  pipe_b_288_0 = _RAND_1088[7:0];
  _RAND_1089 = {1{`RANDOM}};
  pipe_b_288_1 = _RAND_1089[7:0];
  _RAND_1090 = {1{`RANDOM}};
  pipe_b_289_0 = _RAND_1090[19:0];
  _RAND_1091 = {1{`RANDOM}};
  pipe_b_289_1 = _RAND_1091[19:0];
  _RAND_1092 = {1{`RANDOM}};
  pipe_b_290_0 = _RAND_1092[19:0];
  _RAND_1093 = {1{`RANDOM}};
  pipe_b_290_1 = _RAND_1093[19:0];
  _RAND_1094 = {1{`RANDOM}};
  pipe_b_291_0 = _RAND_1094[19:0];
  _RAND_1095 = {1{`RANDOM}};
  pipe_b_291_1 = _RAND_1095[19:0];
  _RAND_1096 = {1{`RANDOM}};
  pipe_b_292_0 = _RAND_1096[19:0];
  _RAND_1097 = {1{`RANDOM}};
  pipe_b_292_1 = _RAND_1097[19:0];
  _RAND_1098 = {1{`RANDOM}};
  pipe_b_293_0 = _RAND_1098[19:0];
  _RAND_1099 = {1{`RANDOM}};
  pipe_b_293_1 = _RAND_1099[19:0];
  _RAND_1100 = {1{`RANDOM}};
  pipe_b_294_0 = _RAND_1100[19:0];
  _RAND_1101 = {1{`RANDOM}};
  pipe_b_294_1 = _RAND_1101[19:0];
  _RAND_1102 = {1{`RANDOM}};
  pipe_b_295_0 = _RAND_1102[19:0];
  _RAND_1103 = {1{`RANDOM}};
  pipe_b_295_1 = _RAND_1103[19:0];
  _RAND_1104 = {1{`RANDOM}};
  pipe_b_296_0 = _RAND_1104[19:0];
  _RAND_1105 = {1{`RANDOM}};
  pipe_b_296_1 = _RAND_1105[19:0];
  _RAND_1106 = {1{`RANDOM}};
  pipe_b_297_0 = _RAND_1106[19:0];
  _RAND_1107 = {1{`RANDOM}};
  pipe_b_297_1 = _RAND_1107[19:0];
  _RAND_1108 = {1{`RANDOM}};
  pipe_b_298_0 = _RAND_1108[19:0];
  _RAND_1109 = {1{`RANDOM}};
  pipe_b_298_1 = _RAND_1109[19:0];
  _RAND_1110 = {1{`RANDOM}};
  pipe_b_299_0 = _RAND_1110[19:0];
  _RAND_1111 = {1{`RANDOM}};
  pipe_b_299_1 = _RAND_1111[19:0];
  _RAND_1112 = {1{`RANDOM}};
  pipe_b_300_0 = _RAND_1112[19:0];
  _RAND_1113 = {1{`RANDOM}};
  pipe_b_300_1 = _RAND_1113[19:0];
  _RAND_1114 = {1{`RANDOM}};
  pipe_b_301_0 = _RAND_1114[19:0];
  _RAND_1115 = {1{`RANDOM}};
  pipe_b_301_1 = _RAND_1115[19:0];
  _RAND_1116 = {1{`RANDOM}};
  pipe_b_302_0 = _RAND_1116[19:0];
  _RAND_1117 = {1{`RANDOM}};
  pipe_b_302_1 = _RAND_1117[19:0];
  _RAND_1118 = {1{`RANDOM}};
  pipe_b_303_0 = _RAND_1118[19:0];
  _RAND_1119 = {1{`RANDOM}};
  pipe_b_303_1 = _RAND_1119[19:0];
  _RAND_1120 = {1{`RANDOM}};
  pipe_b_304_0 = _RAND_1120[7:0];
  _RAND_1121 = {1{`RANDOM}};
  pipe_b_304_1 = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  pipe_b_305_0 = _RAND_1122[19:0];
  _RAND_1123 = {1{`RANDOM}};
  pipe_b_305_1 = _RAND_1123[19:0];
  _RAND_1124 = {1{`RANDOM}};
  pipe_b_306_0 = _RAND_1124[19:0];
  _RAND_1125 = {1{`RANDOM}};
  pipe_b_306_1 = _RAND_1125[19:0];
  _RAND_1126 = {1{`RANDOM}};
  pipe_b_307_0 = _RAND_1126[19:0];
  _RAND_1127 = {1{`RANDOM}};
  pipe_b_307_1 = _RAND_1127[19:0];
  _RAND_1128 = {1{`RANDOM}};
  pipe_b_308_0 = _RAND_1128[19:0];
  _RAND_1129 = {1{`RANDOM}};
  pipe_b_308_1 = _RAND_1129[19:0];
  _RAND_1130 = {1{`RANDOM}};
  pipe_b_309_0 = _RAND_1130[19:0];
  _RAND_1131 = {1{`RANDOM}};
  pipe_b_309_1 = _RAND_1131[19:0];
  _RAND_1132 = {1{`RANDOM}};
  pipe_b_310_0 = _RAND_1132[19:0];
  _RAND_1133 = {1{`RANDOM}};
  pipe_b_310_1 = _RAND_1133[19:0];
  _RAND_1134 = {1{`RANDOM}};
  pipe_b_311_0 = _RAND_1134[19:0];
  _RAND_1135 = {1{`RANDOM}};
  pipe_b_311_1 = _RAND_1135[19:0];
  _RAND_1136 = {1{`RANDOM}};
  pipe_b_312_0 = _RAND_1136[19:0];
  _RAND_1137 = {1{`RANDOM}};
  pipe_b_312_1 = _RAND_1137[19:0];
  _RAND_1138 = {1{`RANDOM}};
  pipe_b_313_0 = _RAND_1138[19:0];
  _RAND_1139 = {1{`RANDOM}};
  pipe_b_313_1 = _RAND_1139[19:0];
  _RAND_1140 = {1{`RANDOM}};
  pipe_b_314_0 = _RAND_1140[19:0];
  _RAND_1141 = {1{`RANDOM}};
  pipe_b_314_1 = _RAND_1141[19:0];
  _RAND_1142 = {1{`RANDOM}};
  pipe_b_315_0 = _RAND_1142[19:0];
  _RAND_1143 = {1{`RANDOM}};
  pipe_b_315_1 = _RAND_1143[19:0];
  _RAND_1144 = {1{`RANDOM}};
  pipe_b_316_0 = _RAND_1144[19:0];
  _RAND_1145 = {1{`RANDOM}};
  pipe_b_316_1 = _RAND_1145[19:0];
  _RAND_1146 = {1{`RANDOM}};
  pipe_b_317_0 = _RAND_1146[19:0];
  _RAND_1147 = {1{`RANDOM}};
  pipe_b_317_1 = _RAND_1147[19:0];
  _RAND_1148 = {1{`RANDOM}};
  pipe_b_318_0 = _RAND_1148[19:0];
  _RAND_1149 = {1{`RANDOM}};
  pipe_b_318_1 = _RAND_1149[19:0];
  _RAND_1150 = {1{`RANDOM}};
  pipe_b_319_0 = _RAND_1150[19:0];
  _RAND_1151 = {1{`RANDOM}};
  pipe_b_319_1 = _RAND_1151[19:0];
  _RAND_1152 = {1{`RANDOM}};
  pipe_b_320_0 = _RAND_1152[7:0];
  _RAND_1153 = {1{`RANDOM}};
  pipe_b_320_1 = _RAND_1153[7:0];
  _RAND_1154 = {1{`RANDOM}};
  pipe_b_321_0 = _RAND_1154[19:0];
  _RAND_1155 = {1{`RANDOM}};
  pipe_b_321_1 = _RAND_1155[19:0];
  _RAND_1156 = {1{`RANDOM}};
  pipe_b_322_0 = _RAND_1156[19:0];
  _RAND_1157 = {1{`RANDOM}};
  pipe_b_322_1 = _RAND_1157[19:0];
  _RAND_1158 = {1{`RANDOM}};
  pipe_b_323_0 = _RAND_1158[19:0];
  _RAND_1159 = {1{`RANDOM}};
  pipe_b_323_1 = _RAND_1159[19:0];
  _RAND_1160 = {1{`RANDOM}};
  pipe_b_324_0 = _RAND_1160[19:0];
  _RAND_1161 = {1{`RANDOM}};
  pipe_b_324_1 = _RAND_1161[19:0];
  _RAND_1162 = {1{`RANDOM}};
  pipe_b_325_0 = _RAND_1162[19:0];
  _RAND_1163 = {1{`RANDOM}};
  pipe_b_325_1 = _RAND_1163[19:0];
  _RAND_1164 = {1{`RANDOM}};
  pipe_b_326_0 = _RAND_1164[19:0];
  _RAND_1165 = {1{`RANDOM}};
  pipe_b_326_1 = _RAND_1165[19:0];
  _RAND_1166 = {1{`RANDOM}};
  pipe_b_327_0 = _RAND_1166[19:0];
  _RAND_1167 = {1{`RANDOM}};
  pipe_b_327_1 = _RAND_1167[19:0];
  _RAND_1168 = {1{`RANDOM}};
  pipe_b_328_0 = _RAND_1168[19:0];
  _RAND_1169 = {1{`RANDOM}};
  pipe_b_328_1 = _RAND_1169[19:0];
  _RAND_1170 = {1{`RANDOM}};
  pipe_b_329_0 = _RAND_1170[19:0];
  _RAND_1171 = {1{`RANDOM}};
  pipe_b_329_1 = _RAND_1171[19:0];
  _RAND_1172 = {1{`RANDOM}};
  pipe_b_330_0 = _RAND_1172[19:0];
  _RAND_1173 = {1{`RANDOM}};
  pipe_b_330_1 = _RAND_1173[19:0];
  _RAND_1174 = {1{`RANDOM}};
  pipe_b_331_0 = _RAND_1174[19:0];
  _RAND_1175 = {1{`RANDOM}};
  pipe_b_331_1 = _RAND_1175[19:0];
  _RAND_1176 = {1{`RANDOM}};
  pipe_b_332_0 = _RAND_1176[19:0];
  _RAND_1177 = {1{`RANDOM}};
  pipe_b_332_1 = _RAND_1177[19:0];
  _RAND_1178 = {1{`RANDOM}};
  pipe_b_333_0 = _RAND_1178[19:0];
  _RAND_1179 = {1{`RANDOM}};
  pipe_b_333_1 = _RAND_1179[19:0];
  _RAND_1180 = {1{`RANDOM}};
  pipe_b_334_0 = _RAND_1180[19:0];
  _RAND_1181 = {1{`RANDOM}};
  pipe_b_334_1 = _RAND_1181[19:0];
  _RAND_1182 = {1{`RANDOM}};
  pipe_b_335_0 = _RAND_1182[19:0];
  _RAND_1183 = {1{`RANDOM}};
  pipe_b_335_1 = _RAND_1183[19:0];
  _RAND_1184 = {1{`RANDOM}};
  pipe_b_336_0 = _RAND_1184[7:0];
  _RAND_1185 = {1{`RANDOM}};
  pipe_b_336_1 = _RAND_1185[7:0];
  _RAND_1186 = {1{`RANDOM}};
  pipe_b_337_0 = _RAND_1186[19:0];
  _RAND_1187 = {1{`RANDOM}};
  pipe_b_337_1 = _RAND_1187[19:0];
  _RAND_1188 = {1{`RANDOM}};
  pipe_b_338_0 = _RAND_1188[19:0];
  _RAND_1189 = {1{`RANDOM}};
  pipe_b_338_1 = _RAND_1189[19:0];
  _RAND_1190 = {1{`RANDOM}};
  pipe_b_339_0 = _RAND_1190[19:0];
  _RAND_1191 = {1{`RANDOM}};
  pipe_b_339_1 = _RAND_1191[19:0];
  _RAND_1192 = {1{`RANDOM}};
  pipe_b_340_0 = _RAND_1192[19:0];
  _RAND_1193 = {1{`RANDOM}};
  pipe_b_340_1 = _RAND_1193[19:0];
  _RAND_1194 = {1{`RANDOM}};
  pipe_b_341_0 = _RAND_1194[19:0];
  _RAND_1195 = {1{`RANDOM}};
  pipe_b_341_1 = _RAND_1195[19:0];
  _RAND_1196 = {1{`RANDOM}};
  pipe_b_342_0 = _RAND_1196[19:0];
  _RAND_1197 = {1{`RANDOM}};
  pipe_b_342_1 = _RAND_1197[19:0];
  _RAND_1198 = {1{`RANDOM}};
  pipe_b_343_0 = _RAND_1198[19:0];
  _RAND_1199 = {1{`RANDOM}};
  pipe_b_343_1 = _RAND_1199[19:0];
  _RAND_1200 = {1{`RANDOM}};
  pipe_b_344_0 = _RAND_1200[19:0];
  _RAND_1201 = {1{`RANDOM}};
  pipe_b_344_1 = _RAND_1201[19:0];
  _RAND_1202 = {1{`RANDOM}};
  pipe_b_345_0 = _RAND_1202[19:0];
  _RAND_1203 = {1{`RANDOM}};
  pipe_b_345_1 = _RAND_1203[19:0];
  _RAND_1204 = {1{`RANDOM}};
  pipe_b_346_0 = _RAND_1204[19:0];
  _RAND_1205 = {1{`RANDOM}};
  pipe_b_346_1 = _RAND_1205[19:0];
  _RAND_1206 = {1{`RANDOM}};
  pipe_b_347_0 = _RAND_1206[19:0];
  _RAND_1207 = {1{`RANDOM}};
  pipe_b_347_1 = _RAND_1207[19:0];
  _RAND_1208 = {1{`RANDOM}};
  pipe_b_348_0 = _RAND_1208[19:0];
  _RAND_1209 = {1{`RANDOM}};
  pipe_b_348_1 = _RAND_1209[19:0];
  _RAND_1210 = {1{`RANDOM}};
  pipe_b_349_0 = _RAND_1210[19:0];
  _RAND_1211 = {1{`RANDOM}};
  pipe_b_349_1 = _RAND_1211[19:0];
  _RAND_1212 = {1{`RANDOM}};
  pipe_b_350_0 = _RAND_1212[19:0];
  _RAND_1213 = {1{`RANDOM}};
  pipe_b_350_1 = _RAND_1213[19:0];
  _RAND_1214 = {1{`RANDOM}};
  pipe_b_351_0 = _RAND_1214[19:0];
  _RAND_1215 = {1{`RANDOM}};
  pipe_b_351_1 = _RAND_1215[19:0];
  _RAND_1216 = {1{`RANDOM}};
  pipe_b_352_0 = _RAND_1216[7:0];
  _RAND_1217 = {1{`RANDOM}};
  pipe_b_352_1 = _RAND_1217[7:0];
  _RAND_1218 = {1{`RANDOM}};
  pipe_b_353_0 = _RAND_1218[19:0];
  _RAND_1219 = {1{`RANDOM}};
  pipe_b_353_1 = _RAND_1219[19:0];
  _RAND_1220 = {1{`RANDOM}};
  pipe_b_354_0 = _RAND_1220[19:0];
  _RAND_1221 = {1{`RANDOM}};
  pipe_b_354_1 = _RAND_1221[19:0];
  _RAND_1222 = {1{`RANDOM}};
  pipe_b_355_0 = _RAND_1222[19:0];
  _RAND_1223 = {1{`RANDOM}};
  pipe_b_355_1 = _RAND_1223[19:0];
  _RAND_1224 = {1{`RANDOM}};
  pipe_b_356_0 = _RAND_1224[19:0];
  _RAND_1225 = {1{`RANDOM}};
  pipe_b_356_1 = _RAND_1225[19:0];
  _RAND_1226 = {1{`RANDOM}};
  pipe_b_357_0 = _RAND_1226[19:0];
  _RAND_1227 = {1{`RANDOM}};
  pipe_b_357_1 = _RAND_1227[19:0];
  _RAND_1228 = {1{`RANDOM}};
  pipe_b_358_0 = _RAND_1228[19:0];
  _RAND_1229 = {1{`RANDOM}};
  pipe_b_358_1 = _RAND_1229[19:0];
  _RAND_1230 = {1{`RANDOM}};
  pipe_b_359_0 = _RAND_1230[19:0];
  _RAND_1231 = {1{`RANDOM}};
  pipe_b_359_1 = _RAND_1231[19:0];
  _RAND_1232 = {1{`RANDOM}};
  pipe_b_360_0 = _RAND_1232[19:0];
  _RAND_1233 = {1{`RANDOM}};
  pipe_b_360_1 = _RAND_1233[19:0];
  _RAND_1234 = {1{`RANDOM}};
  pipe_b_361_0 = _RAND_1234[19:0];
  _RAND_1235 = {1{`RANDOM}};
  pipe_b_361_1 = _RAND_1235[19:0];
  _RAND_1236 = {1{`RANDOM}};
  pipe_b_362_0 = _RAND_1236[19:0];
  _RAND_1237 = {1{`RANDOM}};
  pipe_b_362_1 = _RAND_1237[19:0];
  _RAND_1238 = {1{`RANDOM}};
  pipe_b_363_0 = _RAND_1238[19:0];
  _RAND_1239 = {1{`RANDOM}};
  pipe_b_363_1 = _RAND_1239[19:0];
  _RAND_1240 = {1{`RANDOM}};
  pipe_b_364_0 = _RAND_1240[19:0];
  _RAND_1241 = {1{`RANDOM}};
  pipe_b_364_1 = _RAND_1241[19:0];
  _RAND_1242 = {1{`RANDOM}};
  pipe_b_365_0 = _RAND_1242[19:0];
  _RAND_1243 = {1{`RANDOM}};
  pipe_b_365_1 = _RAND_1243[19:0];
  _RAND_1244 = {1{`RANDOM}};
  pipe_b_366_0 = _RAND_1244[19:0];
  _RAND_1245 = {1{`RANDOM}};
  pipe_b_366_1 = _RAND_1245[19:0];
  _RAND_1246 = {1{`RANDOM}};
  pipe_b_367_0 = _RAND_1246[19:0];
  _RAND_1247 = {1{`RANDOM}};
  pipe_b_367_1 = _RAND_1247[19:0];
  _RAND_1248 = {1{`RANDOM}};
  pipe_b_368_0 = _RAND_1248[7:0];
  _RAND_1249 = {1{`RANDOM}};
  pipe_b_368_1 = _RAND_1249[7:0];
  _RAND_1250 = {1{`RANDOM}};
  pipe_b_369_0 = _RAND_1250[19:0];
  _RAND_1251 = {1{`RANDOM}};
  pipe_b_369_1 = _RAND_1251[19:0];
  _RAND_1252 = {1{`RANDOM}};
  pipe_b_370_0 = _RAND_1252[19:0];
  _RAND_1253 = {1{`RANDOM}};
  pipe_b_370_1 = _RAND_1253[19:0];
  _RAND_1254 = {1{`RANDOM}};
  pipe_b_371_0 = _RAND_1254[19:0];
  _RAND_1255 = {1{`RANDOM}};
  pipe_b_371_1 = _RAND_1255[19:0];
  _RAND_1256 = {1{`RANDOM}};
  pipe_b_372_0 = _RAND_1256[19:0];
  _RAND_1257 = {1{`RANDOM}};
  pipe_b_372_1 = _RAND_1257[19:0];
  _RAND_1258 = {1{`RANDOM}};
  pipe_b_373_0 = _RAND_1258[19:0];
  _RAND_1259 = {1{`RANDOM}};
  pipe_b_373_1 = _RAND_1259[19:0];
  _RAND_1260 = {1{`RANDOM}};
  pipe_b_374_0 = _RAND_1260[19:0];
  _RAND_1261 = {1{`RANDOM}};
  pipe_b_374_1 = _RAND_1261[19:0];
  _RAND_1262 = {1{`RANDOM}};
  pipe_b_375_0 = _RAND_1262[19:0];
  _RAND_1263 = {1{`RANDOM}};
  pipe_b_375_1 = _RAND_1263[19:0];
  _RAND_1264 = {1{`RANDOM}};
  pipe_b_376_0 = _RAND_1264[19:0];
  _RAND_1265 = {1{`RANDOM}};
  pipe_b_376_1 = _RAND_1265[19:0];
  _RAND_1266 = {1{`RANDOM}};
  pipe_b_377_0 = _RAND_1266[19:0];
  _RAND_1267 = {1{`RANDOM}};
  pipe_b_377_1 = _RAND_1267[19:0];
  _RAND_1268 = {1{`RANDOM}};
  pipe_b_378_0 = _RAND_1268[19:0];
  _RAND_1269 = {1{`RANDOM}};
  pipe_b_378_1 = _RAND_1269[19:0];
  _RAND_1270 = {1{`RANDOM}};
  pipe_b_379_0 = _RAND_1270[19:0];
  _RAND_1271 = {1{`RANDOM}};
  pipe_b_379_1 = _RAND_1271[19:0];
  _RAND_1272 = {1{`RANDOM}};
  pipe_b_380_0 = _RAND_1272[19:0];
  _RAND_1273 = {1{`RANDOM}};
  pipe_b_380_1 = _RAND_1273[19:0];
  _RAND_1274 = {1{`RANDOM}};
  pipe_b_381_0 = _RAND_1274[19:0];
  _RAND_1275 = {1{`RANDOM}};
  pipe_b_381_1 = _RAND_1275[19:0];
  _RAND_1276 = {1{`RANDOM}};
  pipe_b_382_0 = _RAND_1276[19:0];
  _RAND_1277 = {1{`RANDOM}};
  pipe_b_382_1 = _RAND_1277[19:0];
  _RAND_1278 = {1{`RANDOM}};
  pipe_b_383_0 = _RAND_1278[19:0];
  _RAND_1279 = {1{`RANDOM}};
  pipe_b_383_1 = _RAND_1279[19:0];
  _RAND_1280 = {1{`RANDOM}};
  pipe_b_384_0 = _RAND_1280[7:0];
  _RAND_1281 = {1{`RANDOM}};
  pipe_b_384_1 = _RAND_1281[7:0];
  _RAND_1282 = {1{`RANDOM}};
  pipe_b_385_0 = _RAND_1282[19:0];
  _RAND_1283 = {1{`RANDOM}};
  pipe_b_385_1 = _RAND_1283[19:0];
  _RAND_1284 = {1{`RANDOM}};
  pipe_b_386_0 = _RAND_1284[19:0];
  _RAND_1285 = {1{`RANDOM}};
  pipe_b_386_1 = _RAND_1285[19:0];
  _RAND_1286 = {1{`RANDOM}};
  pipe_b_387_0 = _RAND_1286[19:0];
  _RAND_1287 = {1{`RANDOM}};
  pipe_b_387_1 = _RAND_1287[19:0];
  _RAND_1288 = {1{`RANDOM}};
  pipe_b_388_0 = _RAND_1288[19:0];
  _RAND_1289 = {1{`RANDOM}};
  pipe_b_388_1 = _RAND_1289[19:0];
  _RAND_1290 = {1{`RANDOM}};
  pipe_b_389_0 = _RAND_1290[19:0];
  _RAND_1291 = {1{`RANDOM}};
  pipe_b_389_1 = _RAND_1291[19:0];
  _RAND_1292 = {1{`RANDOM}};
  pipe_b_390_0 = _RAND_1292[19:0];
  _RAND_1293 = {1{`RANDOM}};
  pipe_b_390_1 = _RAND_1293[19:0];
  _RAND_1294 = {1{`RANDOM}};
  pipe_b_391_0 = _RAND_1294[19:0];
  _RAND_1295 = {1{`RANDOM}};
  pipe_b_391_1 = _RAND_1295[19:0];
  _RAND_1296 = {1{`RANDOM}};
  pipe_b_392_0 = _RAND_1296[19:0];
  _RAND_1297 = {1{`RANDOM}};
  pipe_b_392_1 = _RAND_1297[19:0];
  _RAND_1298 = {1{`RANDOM}};
  pipe_b_393_0 = _RAND_1298[19:0];
  _RAND_1299 = {1{`RANDOM}};
  pipe_b_393_1 = _RAND_1299[19:0];
  _RAND_1300 = {1{`RANDOM}};
  pipe_b_394_0 = _RAND_1300[19:0];
  _RAND_1301 = {1{`RANDOM}};
  pipe_b_394_1 = _RAND_1301[19:0];
  _RAND_1302 = {1{`RANDOM}};
  pipe_b_395_0 = _RAND_1302[19:0];
  _RAND_1303 = {1{`RANDOM}};
  pipe_b_395_1 = _RAND_1303[19:0];
  _RAND_1304 = {1{`RANDOM}};
  pipe_b_396_0 = _RAND_1304[19:0];
  _RAND_1305 = {1{`RANDOM}};
  pipe_b_396_1 = _RAND_1305[19:0];
  _RAND_1306 = {1{`RANDOM}};
  pipe_b_397_0 = _RAND_1306[19:0];
  _RAND_1307 = {1{`RANDOM}};
  pipe_b_397_1 = _RAND_1307[19:0];
  _RAND_1308 = {1{`RANDOM}};
  pipe_b_398_0 = _RAND_1308[19:0];
  _RAND_1309 = {1{`RANDOM}};
  pipe_b_398_1 = _RAND_1309[19:0];
  _RAND_1310 = {1{`RANDOM}};
  pipe_b_399_0 = _RAND_1310[19:0];
  _RAND_1311 = {1{`RANDOM}};
  pipe_b_399_1 = _RAND_1311[19:0];
  _RAND_1312 = {1{`RANDOM}};
  pipe_b_400_0 = _RAND_1312[7:0];
  _RAND_1313 = {1{`RANDOM}};
  pipe_b_400_1 = _RAND_1313[7:0];
  _RAND_1314 = {1{`RANDOM}};
  pipe_b_401_0 = _RAND_1314[19:0];
  _RAND_1315 = {1{`RANDOM}};
  pipe_b_401_1 = _RAND_1315[19:0];
  _RAND_1316 = {1{`RANDOM}};
  pipe_b_402_0 = _RAND_1316[19:0];
  _RAND_1317 = {1{`RANDOM}};
  pipe_b_402_1 = _RAND_1317[19:0];
  _RAND_1318 = {1{`RANDOM}};
  pipe_b_403_0 = _RAND_1318[19:0];
  _RAND_1319 = {1{`RANDOM}};
  pipe_b_403_1 = _RAND_1319[19:0];
  _RAND_1320 = {1{`RANDOM}};
  pipe_b_404_0 = _RAND_1320[19:0];
  _RAND_1321 = {1{`RANDOM}};
  pipe_b_404_1 = _RAND_1321[19:0];
  _RAND_1322 = {1{`RANDOM}};
  pipe_b_405_0 = _RAND_1322[19:0];
  _RAND_1323 = {1{`RANDOM}};
  pipe_b_405_1 = _RAND_1323[19:0];
  _RAND_1324 = {1{`RANDOM}};
  pipe_b_406_0 = _RAND_1324[19:0];
  _RAND_1325 = {1{`RANDOM}};
  pipe_b_406_1 = _RAND_1325[19:0];
  _RAND_1326 = {1{`RANDOM}};
  pipe_b_407_0 = _RAND_1326[19:0];
  _RAND_1327 = {1{`RANDOM}};
  pipe_b_407_1 = _RAND_1327[19:0];
  _RAND_1328 = {1{`RANDOM}};
  pipe_b_408_0 = _RAND_1328[19:0];
  _RAND_1329 = {1{`RANDOM}};
  pipe_b_408_1 = _RAND_1329[19:0];
  _RAND_1330 = {1{`RANDOM}};
  pipe_b_409_0 = _RAND_1330[19:0];
  _RAND_1331 = {1{`RANDOM}};
  pipe_b_409_1 = _RAND_1331[19:0];
  _RAND_1332 = {1{`RANDOM}};
  pipe_b_410_0 = _RAND_1332[19:0];
  _RAND_1333 = {1{`RANDOM}};
  pipe_b_410_1 = _RAND_1333[19:0];
  _RAND_1334 = {1{`RANDOM}};
  pipe_b_411_0 = _RAND_1334[19:0];
  _RAND_1335 = {1{`RANDOM}};
  pipe_b_411_1 = _RAND_1335[19:0];
  _RAND_1336 = {1{`RANDOM}};
  pipe_b_412_0 = _RAND_1336[19:0];
  _RAND_1337 = {1{`RANDOM}};
  pipe_b_412_1 = _RAND_1337[19:0];
  _RAND_1338 = {1{`RANDOM}};
  pipe_b_413_0 = _RAND_1338[19:0];
  _RAND_1339 = {1{`RANDOM}};
  pipe_b_413_1 = _RAND_1339[19:0];
  _RAND_1340 = {1{`RANDOM}};
  pipe_b_414_0 = _RAND_1340[19:0];
  _RAND_1341 = {1{`RANDOM}};
  pipe_b_414_1 = _RAND_1341[19:0];
  _RAND_1342 = {1{`RANDOM}};
  pipe_b_415_0 = _RAND_1342[19:0];
  _RAND_1343 = {1{`RANDOM}};
  pipe_b_415_1 = _RAND_1343[19:0];
  _RAND_1344 = {1{`RANDOM}};
  pipe_b_416_0 = _RAND_1344[7:0];
  _RAND_1345 = {1{`RANDOM}};
  pipe_b_416_1 = _RAND_1345[7:0];
  _RAND_1346 = {1{`RANDOM}};
  pipe_b_417_0 = _RAND_1346[19:0];
  _RAND_1347 = {1{`RANDOM}};
  pipe_b_417_1 = _RAND_1347[19:0];
  _RAND_1348 = {1{`RANDOM}};
  pipe_b_418_0 = _RAND_1348[19:0];
  _RAND_1349 = {1{`RANDOM}};
  pipe_b_418_1 = _RAND_1349[19:0];
  _RAND_1350 = {1{`RANDOM}};
  pipe_b_419_0 = _RAND_1350[19:0];
  _RAND_1351 = {1{`RANDOM}};
  pipe_b_419_1 = _RAND_1351[19:0];
  _RAND_1352 = {1{`RANDOM}};
  pipe_b_420_0 = _RAND_1352[19:0];
  _RAND_1353 = {1{`RANDOM}};
  pipe_b_420_1 = _RAND_1353[19:0];
  _RAND_1354 = {1{`RANDOM}};
  pipe_b_421_0 = _RAND_1354[19:0];
  _RAND_1355 = {1{`RANDOM}};
  pipe_b_421_1 = _RAND_1355[19:0];
  _RAND_1356 = {1{`RANDOM}};
  pipe_b_422_0 = _RAND_1356[19:0];
  _RAND_1357 = {1{`RANDOM}};
  pipe_b_422_1 = _RAND_1357[19:0];
  _RAND_1358 = {1{`RANDOM}};
  pipe_b_423_0 = _RAND_1358[19:0];
  _RAND_1359 = {1{`RANDOM}};
  pipe_b_423_1 = _RAND_1359[19:0];
  _RAND_1360 = {1{`RANDOM}};
  pipe_b_424_0 = _RAND_1360[19:0];
  _RAND_1361 = {1{`RANDOM}};
  pipe_b_424_1 = _RAND_1361[19:0];
  _RAND_1362 = {1{`RANDOM}};
  pipe_b_425_0 = _RAND_1362[19:0];
  _RAND_1363 = {1{`RANDOM}};
  pipe_b_425_1 = _RAND_1363[19:0];
  _RAND_1364 = {1{`RANDOM}};
  pipe_b_426_0 = _RAND_1364[19:0];
  _RAND_1365 = {1{`RANDOM}};
  pipe_b_426_1 = _RAND_1365[19:0];
  _RAND_1366 = {1{`RANDOM}};
  pipe_b_427_0 = _RAND_1366[19:0];
  _RAND_1367 = {1{`RANDOM}};
  pipe_b_427_1 = _RAND_1367[19:0];
  _RAND_1368 = {1{`RANDOM}};
  pipe_b_428_0 = _RAND_1368[19:0];
  _RAND_1369 = {1{`RANDOM}};
  pipe_b_428_1 = _RAND_1369[19:0];
  _RAND_1370 = {1{`RANDOM}};
  pipe_b_429_0 = _RAND_1370[19:0];
  _RAND_1371 = {1{`RANDOM}};
  pipe_b_429_1 = _RAND_1371[19:0];
  _RAND_1372 = {1{`RANDOM}};
  pipe_b_430_0 = _RAND_1372[19:0];
  _RAND_1373 = {1{`RANDOM}};
  pipe_b_430_1 = _RAND_1373[19:0];
  _RAND_1374 = {1{`RANDOM}};
  pipe_b_431_0 = _RAND_1374[19:0];
  _RAND_1375 = {1{`RANDOM}};
  pipe_b_431_1 = _RAND_1375[19:0];
  _RAND_1376 = {1{`RANDOM}};
  pipe_b_432_0 = _RAND_1376[7:0];
  _RAND_1377 = {1{`RANDOM}};
  pipe_b_432_1 = _RAND_1377[7:0];
  _RAND_1378 = {1{`RANDOM}};
  pipe_b_433_0 = _RAND_1378[19:0];
  _RAND_1379 = {1{`RANDOM}};
  pipe_b_433_1 = _RAND_1379[19:0];
  _RAND_1380 = {1{`RANDOM}};
  pipe_b_434_0 = _RAND_1380[19:0];
  _RAND_1381 = {1{`RANDOM}};
  pipe_b_434_1 = _RAND_1381[19:0];
  _RAND_1382 = {1{`RANDOM}};
  pipe_b_435_0 = _RAND_1382[19:0];
  _RAND_1383 = {1{`RANDOM}};
  pipe_b_435_1 = _RAND_1383[19:0];
  _RAND_1384 = {1{`RANDOM}};
  pipe_b_436_0 = _RAND_1384[19:0];
  _RAND_1385 = {1{`RANDOM}};
  pipe_b_436_1 = _RAND_1385[19:0];
  _RAND_1386 = {1{`RANDOM}};
  pipe_b_437_0 = _RAND_1386[19:0];
  _RAND_1387 = {1{`RANDOM}};
  pipe_b_437_1 = _RAND_1387[19:0];
  _RAND_1388 = {1{`RANDOM}};
  pipe_b_438_0 = _RAND_1388[19:0];
  _RAND_1389 = {1{`RANDOM}};
  pipe_b_438_1 = _RAND_1389[19:0];
  _RAND_1390 = {1{`RANDOM}};
  pipe_b_439_0 = _RAND_1390[19:0];
  _RAND_1391 = {1{`RANDOM}};
  pipe_b_439_1 = _RAND_1391[19:0];
  _RAND_1392 = {1{`RANDOM}};
  pipe_b_440_0 = _RAND_1392[19:0];
  _RAND_1393 = {1{`RANDOM}};
  pipe_b_440_1 = _RAND_1393[19:0];
  _RAND_1394 = {1{`RANDOM}};
  pipe_b_441_0 = _RAND_1394[19:0];
  _RAND_1395 = {1{`RANDOM}};
  pipe_b_441_1 = _RAND_1395[19:0];
  _RAND_1396 = {1{`RANDOM}};
  pipe_b_442_0 = _RAND_1396[19:0];
  _RAND_1397 = {1{`RANDOM}};
  pipe_b_442_1 = _RAND_1397[19:0];
  _RAND_1398 = {1{`RANDOM}};
  pipe_b_443_0 = _RAND_1398[19:0];
  _RAND_1399 = {1{`RANDOM}};
  pipe_b_443_1 = _RAND_1399[19:0];
  _RAND_1400 = {1{`RANDOM}};
  pipe_b_444_0 = _RAND_1400[19:0];
  _RAND_1401 = {1{`RANDOM}};
  pipe_b_444_1 = _RAND_1401[19:0];
  _RAND_1402 = {1{`RANDOM}};
  pipe_b_445_0 = _RAND_1402[19:0];
  _RAND_1403 = {1{`RANDOM}};
  pipe_b_445_1 = _RAND_1403[19:0];
  _RAND_1404 = {1{`RANDOM}};
  pipe_b_446_0 = _RAND_1404[19:0];
  _RAND_1405 = {1{`RANDOM}};
  pipe_b_446_1 = _RAND_1405[19:0];
  _RAND_1406 = {1{`RANDOM}};
  pipe_b_447_0 = _RAND_1406[19:0];
  _RAND_1407 = {1{`RANDOM}};
  pipe_b_447_1 = _RAND_1407[19:0];
  _RAND_1408 = {1{`RANDOM}};
  pipe_b_448_0 = _RAND_1408[7:0];
  _RAND_1409 = {1{`RANDOM}};
  pipe_b_448_1 = _RAND_1409[7:0];
  _RAND_1410 = {1{`RANDOM}};
  pipe_b_449_0 = _RAND_1410[19:0];
  _RAND_1411 = {1{`RANDOM}};
  pipe_b_449_1 = _RAND_1411[19:0];
  _RAND_1412 = {1{`RANDOM}};
  pipe_b_450_0 = _RAND_1412[19:0];
  _RAND_1413 = {1{`RANDOM}};
  pipe_b_450_1 = _RAND_1413[19:0];
  _RAND_1414 = {1{`RANDOM}};
  pipe_b_451_0 = _RAND_1414[19:0];
  _RAND_1415 = {1{`RANDOM}};
  pipe_b_451_1 = _RAND_1415[19:0];
  _RAND_1416 = {1{`RANDOM}};
  pipe_b_452_0 = _RAND_1416[19:0];
  _RAND_1417 = {1{`RANDOM}};
  pipe_b_452_1 = _RAND_1417[19:0];
  _RAND_1418 = {1{`RANDOM}};
  pipe_b_453_0 = _RAND_1418[19:0];
  _RAND_1419 = {1{`RANDOM}};
  pipe_b_453_1 = _RAND_1419[19:0];
  _RAND_1420 = {1{`RANDOM}};
  pipe_b_454_0 = _RAND_1420[19:0];
  _RAND_1421 = {1{`RANDOM}};
  pipe_b_454_1 = _RAND_1421[19:0];
  _RAND_1422 = {1{`RANDOM}};
  pipe_b_455_0 = _RAND_1422[19:0];
  _RAND_1423 = {1{`RANDOM}};
  pipe_b_455_1 = _RAND_1423[19:0];
  _RAND_1424 = {1{`RANDOM}};
  pipe_b_456_0 = _RAND_1424[19:0];
  _RAND_1425 = {1{`RANDOM}};
  pipe_b_456_1 = _RAND_1425[19:0];
  _RAND_1426 = {1{`RANDOM}};
  pipe_b_457_0 = _RAND_1426[19:0];
  _RAND_1427 = {1{`RANDOM}};
  pipe_b_457_1 = _RAND_1427[19:0];
  _RAND_1428 = {1{`RANDOM}};
  pipe_b_458_0 = _RAND_1428[19:0];
  _RAND_1429 = {1{`RANDOM}};
  pipe_b_458_1 = _RAND_1429[19:0];
  _RAND_1430 = {1{`RANDOM}};
  pipe_b_459_0 = _RAND_1430[19:0];
  _RAND_1431 = {1{`RANDOM}};
  pipe_b_459_1 = _RAND_1431[19:0];
  _RAND_1432 = {1{`RANDOM}};
  pipe_b_460_0 = _RAND_1432[19:0];
  _RAND_1433 = {1{`RANDOM}};
  pipe_b_460_1 = _RAND_1433[19:0];
  _RAND_1434 = {1{`RANDOM}};
  pipe_b_461_0 = _RAND_1434[19:0];
  _RAND_1435 = {1{`RANDOM}};
  pipe_b_461_1 = _RAND_1435[19:0];
  _RAND_1436 = {1{`RANDOM}};
  pipe_b_462_0 = _RAND_1436[19:0];
  _RAND_1437 = {1{`RANDOM}};
  pipe_b_462_1 = _RAND_1437[19:0];
  _RAND_1438 = {1{`RANDOM}};
  pipe_b_463_0 = _RAND_1438[19:0];
  _RAND_1439 = {1{`RANDOM}};
  pipe_b_463_1 = _RAND_1439[19:0];
  _RAND_1440 = {1{`RANDOM}};
  pipe_b_464_0 = _RAND_1440[7:0];
  _RAND_1441 = {1{`RANDOM}};
  pipe_b_464_1 = _RAND_1441[7:0];
  _RAND_1442 = {1{`RANDOM}};
  pipe_b_465_0 = _RAND_1442[19:0];
  _RAND_1443 = {1{`RANDOM}};
  pipe_b_465_1 = _RAND_1443[19:0];
  _RAND_1444 = {1{`RANDOM}};
  pipe_b_466_0 = _RAND_1444[19:0];
  _RAND_1445 = {1{`RANDOM}};
  pipe_b_466_1 = _RAND_1445[19:0];
  _RAND_1446 = {1{`RANDOM}};
  pipe_b_467_0 = _RAND_1446[19:0];
  _RAND_1447 = {1{`RANDOM}};
  pipe_b_467_1 = _RAND_1447[19:0];
  _RAND_1448 = {1{`RANDOM}};
  pipe_b_468_0 = _RAND_1448[19:0];
  _RAND_1449 = {1{`RANDOM}};
  pipe_b_468_1 = _RAND_1449[19:0];
  _RAND_1450 = {1{`RANDOM}};
  pipe_b_469_0 = _RAND_1450[19:0];
  _RAND_1451 = {1{`RANDOM}};
  pipe_b_469_1 = _RAND_1451[19:0];
  _RAND_1452 = {1{`RANDOM}};
  pipe_b_470_0 = _RAND_1452[19:0];
  _RAND_1453 = {1{`RANDOM}};
  pipe_b_470_1 = _RAND_1453[19:0];
  _RAND_1454 = {1{`RANDOM}};
  pipe_b_471_0 = _RAND_1454[19:0];
  _RAND_1455 = {1{`RANDOM}};
  pipe_b_471_1 = _RAND_1455[19:0];
  _RAND_1456 = {1{`RANDOM}};
  pipe_b_472_0 = _RAND_1456[19:0];
  _RAND_1457 = {1{`RANDOM}};
  pipe_b_472_1 = _RAND_1457[19:0];
  _RAND_1458 = {1{`RANDOM}};
  pipe_b_473_0 = _RAND_1458[19:0];
  _RAND_1459 = {1{`RANDOM}};
  pipe_b_473_1 = _RAND_1459[19:0];
  _RAND_1460 = {1{`RANDOM}};
  pipe_b_474_0 = _RAND_1460[19:0];
  _RAND_1461 = {1{`RANDOM}};
  pipe_b_474_1 = _RAND_1461[19:0];
  _RAND_1462 = {1{`RANDOM}};
  pipe_b_475_0 = _RAND_1462[19:0];
  _RAND_1463 = {1{`RANDOM}};
  pipe_b_475_1 = _RAND_1463[19:0];
  _RAND_1464 = {1{`RANDOM}};
  pipe_b_476_0 = _RAND_1464[19:0];
  _RAND_1465 = {1{`RANDOM}};
  pipe_b_476_1 = _RAND_1465[19:0];
  _RAND_1466 = {1{`RANDOM}};
  pipe_b_477_0 = _RAND_1466[19:0];
  _RAND_1467 = {1{`RANDOM}};
  pipe_b_477_1 = _RAND_1467[19:0];
  _RAND_1468 = {1{`RANDOM}};
  pipe_b_478_0 = _RAND_1468[19:0];
  _RAND_1469 = {1{`RANDOM}};
  pipe_b_478_1 = _RAND_1469[19:0];
  _RAND_1470 = {1{`RANDOM}};
  pipe_b_479_0 = _RAND_1470[19:0];
  _RAND_1471 = {1{`RANDOM}};
  pipe_b_479_1 = _RAND_1471[19:0];
  _RAND_1472 = {1{`RANDOM}};
  pipe_b_480_0 = _RAND_1472[7:0];
  _RAND_1473 = {1{`RANDOM}};
  pipe_b_480_1 = _RAND_1473[7:0];
  _RAND_1474 = {1{`RANDOM}};
  pipe_b_481_0 = _RAND_1474[19:0];
  _RAND_1475 = {1{`RANDOM}};
  pipe_b_481_1 = _RAND_1475[19:0];
  _RAND_1476 = {1{`RANDOM}};
  pipe_b_482_0 = _RAND_1476[19:0];
  _RAND_1477 = {1{`RANDOM}};
  pipe_b_482_1 = _RAND_1477[19:0];
  _RAND_1478 = {1{`RANDOM}};
  pipe_b_483_0 = _RAND_1478[19:0];
  _RAND_1479 = {1{`RANDOM}};
  pipe_b_483_1 = _RAND_1479[19:0];
  _RAND_1480 = {1{`RANDOM}};
  pipe_b_484_0 = _RAND_1480[19:0];
  _RAND_1481 = {1{`RANDOM}};
  pipe_b_484_1 = _RAND_1481[19:0];
  _RAND_1482 = {1{`RANDOM}};
  pipe_b_485_0 = _RAND_1482[19:0];
  _RAND_1483 = {1{`RANDOM}};
  pipe_b_485_1 = _RAND_1483[19:0];
  _RAND_1484 = {1{`RANDOM}};
  pipe_b_486_0 = _RAND_1484[19:0];
  _RAND_1485 = {1{`RANDOM}};
  pipe_b_486_1 = _RAND_1485[19:0];
  _RAND_1486 = {1{`RANDOM}};
  pipe_b_487_0 = _RAND_1486[19:0];
  _RAND_1487 = {1{`RANDOM}};
  pipe_b_487_1 = _RAND_1487[19:0];
  _RAND_1488 = {1{`RANDOM}};
  pipe_b_488_0 = _RAND_1488[19:0];
  _RAND_1489 = {1{`RANDOM}};
  pipe_b_488_1 = _RAND_1489[19:0];
  _RAND_1490 = {1{`RANDOM}};
  pipe_b_489_0 = _RAND_1490[19:0];
  _RAND_1491 = {1{`RANDOM}};
  pipe_b_489_1 = _RAND_1491[19:0];
  _RAND_1492 = {1{`RANDOM}};
  pipe_b_490_0 = _RAND_1492[19:0];
  _RAND_1493 = {1{`RANDOM}};
  pipe_b_490_1 = _RAND_1493[19:0];
  _RAND_1494 = {1{`RANDOM}};
  pipe_b_491_0 = _RAND_1494[19:0];
  _RAND_1495 = {1{`RANDOM}};
  pipe_b_491_1 = _RAND_1495[19:0];
  _RAND_1496 = {1{`RANDOM}};
  pipe_b_492_0 = _RAND_1496[19:0];
  _RAND_1497 = {1{`RANDOM}};
  pipe_b_492_1 = _RAND_1497[19:0];
  _RAND_1498 = {1{`RANDOM}};
  pipe_b_493_0 = _RAND_1498[19:0];
  _RAND_1499 = {1{`RANDOM}};
  pipe_b_493_1 = _RAND_1499[19:0];
  _RAND_1500 = {1{`RANDOM}};
  pipe_b_494_0 = _RAND_1500[19:0];
  _RAND_1501 = {1{`RANDOM}};
  pipe_b_494_1 = _RAND_1501[19:0];
  _RAND_1502 = {1{`RANDOM}};
  pipe_b_495_0 = _RAND_1502[19:0];
  _RAND_1503 = {1{`RANDOM}};
  pipe_b_495_1 = _RAND_1503[19:0];
  _RAND_1504 = {1{`RANDOM}};
  pipe_b_496_0 = _RAND_1504[7:0];
  _RAND_1505 = {1{`RANDOM}};
  pipe_b_496_1 = _RAND_1505[7:0];
  _RAND_1506 = {1{`RANDOM}};
  pipe_b_497_0 = _RAND_1506[19:0];
  _RAND_1507 = {1{`RANDOM}};
  pipe_b_497_1 = _RAND_1507[19:0];
  _RAND_1508 = {1{`RANDOM}};
  pipe_b_498_0 = _RAND_1508[19:0];
  _RAND_1509 = {1{`RANDOM}};
  pipe_b_498_1 = _RAND_1509[19:0];
  _RAND_1510 = {1{`RANDOM}};
  pipe_b_499_0 = _RAND_1510[19:0];
  _RAND_1511 = {1{`RANDOM}};
  pipe_b_499_1 = _RAND_1511[19:0];
  _RAND_1512 = {1{`RANDOM}};
  pipe_b_500_0 = _RAND_1512[19:0];
  _RAND_1513 = {1{`RANDOM}};
  pipe_b_500_1 = _RAND_1513[19:0];
  _RAND_1514 = {1{`RANDOM}};
  pipe_b_501_0 = _RAND_1514[19:0];
  _RAND_1515 = {1{`RANDOM}};
  pipe_b_501_1 = _RAND_1515[19:0];
  _RAND_1516 = {1{`RANDOM}};
  pipe_b_502_0 = _RAND_1516[19:0];
  _RAND_1517 = {1{`RANDOM}};
  pipe_b_502_1 = _RAND_1517[19:0];
  _RAND_1518 = {1{`RANDOM}};
  pipe_b_503_0 = _RAND_1518[19:0];
  _RAND_1519 = {1{`RANDOM}};
  pipe_b_503_1 = _RAND_1519[19:0];
  _RAND_1520 = {1{`RANDOM}};
  pipe_b_504_0 = _RAND_1520[19:0];
  _RAND_1521 = {1{`RANDOM}};
  pipe_b_504_1 = _RAND_1521[19:0];
  _RAND_1522 = {1{`RANDOM}};
  pipe_b_505_0 = _RAND_1522[19:0];
  _RAND_1523 = {1{`RANDOM}};
  pipe_b_505_1 = _RAND_1523[19:0];
  _RAND_1524 = {1{`RANDOM}};
  pipe_b_506_0 = _RAND_1524[19:0];
  _RAND_1525 = {1{`RANDOM}};
  pipe_b_506_1 = _RAND_1525[19:0];
  _RAND_1526 = {1{`RANDOM}};
  pipe_b_507_0 = _RAND_1526[19:0];
  _RAND_1527 = {1{`RANDOM}};
  pipe_b_507_1 = _RAND_1527[19:0];
  _RAND_1528 = {1{`RANDOM}};
  pipe_b_508_0 = _RAND_1528[19:0];
  _RAND_1529 = {1{`RANDOM}};
  pipe_b_508_1 = _RAND_1529[19:0];
  _RAND_1530 = {1{`RANDOM}};
  pipe_b_509_0 = _RAND_1530[19:0];
  _RAND_1531 = {1{`RANDOM}};
  pipe_b_509_1 = _RAND_1531[19:0];
  _RAND_1532 = {1{`RANDOM}};
  pipe_b_510_0 = _RAND_1532[19:0];
  _RAND_1533 = {1{`RANDOM}};
  pipe_b_510_1 = _RAND_1533[19:0];
  _RAND_1534 = {1{`RANDOM}};
  pipe_b_511_0 = _RAND_1534[19:0];
  _RAND_1535 = {1{`RANDOM}};
  pipe_b_511_1 = _RAND_1535[19:0];
  _RAND_1536 = {1{`RANDOM}};
  mesh_0_0_io_in_control_0_shift_pipe_b = _RAND_1536[4:0];
  _RAND_1537 = {1{`RANDOM}};
  mesh_0_0_io_in_control_0_dataflow_pipe_b = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  mesh_0_0_io_in_control_0_propagate_pipe_b = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  mesh_0_0_io_in_control_1_shift_pipe_b = _RAND_1539[4:0];
  _RAND_1540 = {1{`RANDOM}};
  mesh_0_0_io_in_control_1_dataflow_pipe_b = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  mesh_0_0_io_in_control_1_propagate_pipe_b = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  mesh_1_0_io_in_control_0_shift_pipe_b = _RAND_1542[4:0];
  _RAND_1543 = {1{`RANDOM}};
  mesh_1_0_io_in_control_0_dataflow_pipe_b = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  mesh_1_0_io_in_control_0_propagate_pipe_b = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  mesh_1_0_io_in_control_1_shift_pipe_b = _RAND_1545[4:0];
  _RAND_1546 = {1{`RANDOM}};
  mesh_1_0_io_in_control_1_dataflow_pipe_b = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  mesh_1_0_io_in_control_1_propagate_pipe_b = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  mesh_2_0_io_in_control_0_shift_pipe_b = _RAND_1548[4:0];
  _RAND_1549 = {1{`RANDOM}};
  mesh_2_0_io_in_control_0_dataflow_pipe_b = _RAND_1549[0:0];
  _RAND_1550 = {1{`RANDOM}};
  mesh_2_0_io_in_control_0_propagate_pipe_b = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  mesh_2_0_io_in_control_1_shift_pipe_b = _RAND_1551[4:0];
  _RAND_1552 = {1{`RANDOM}};
  mesh_2_0_io_in_control_1_dataflow_pipe_b = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  mesh_2_0_io_in_control_1_propagate_pipe_b = _RAND_1553[0:0];
  _RAND_1554 = {1{`RANDOM}};
  mesh_3_0_io_in_control_0_shift_pipe_b = _RAND_1554[4:0];
  _RAND_1555 = {1{`RANDOM}};
  mesh_3_0_io_in_control_0_dataflow_pipe_b = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  mesh_3_0_io_in_control_0_propagate_pipe_b = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  mesh_3_0_io_in_control_1_shift_pipe_b = _RAND_1557[4:0];
  _RAND_1558 = {1{`RANDOM}};
  mesh_3_0_io_in_control_1_dataflow_pipe_b = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  mesh_3_0_io_in_control_1_propagate_pipe_b = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  mesh_4_0_io_in_control_0_shift_pipe_b = _RAND_1560[4:0];
  _RAND_1561 = {1{`RANDOM}};
  mesh_4_0_io_in_control_0_dataflow_pipe_b = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  mesh_4_0_io_in_control_0_propagate_pipe_b = _RAND_1562[0:0];
  _RAND_1563 = {1{`RANDOM}};
  mesh_4_0_io_in_control_1_shift_pipe_b = _RAND_1563[4:0];
  _RAND_1564 = {1{`RANDOM}};
  mesh_4_0_io_in_control_1_dataflow_pipe_b = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  mesh_4_0_io_in_control_1_propagate_pipe_b = _RAND_1565[0:0];
  _RAND_1566 = {1{`RANDOM}};
  mesh_5_0_io_in_control_0_shift_pipe_b = _RAND_1566[4:0];
  _RAND_1567 = {1{`RANDOM}};
  mesh_5_0_io_in_control_0_dataflow_pipe_b = _RAND_1567[0:0];
  _RAND_1568 = {1{`RANDOM}};
  mesh_5_0_io_in_control_0_propagate_pipe_b = _RAND_1568[0:0];
  _RAND_1569 = {1{`RANDOM}};
  mesh_5_0_io_in_control_1_shift_pipe_b = _RAND_1569[4:0];
  _RAND_1570 = {1{`RANDOM}};
  mesh_5_0_io_in_control_1_dataflow_pipe_b = _RAND_1570[0:0];
  _RAND_1571 = {1{`RANDOM}};
  mesh_5_0_io_in_control_1_propagate_pipe_b = _RAND_1571[0:0];
  _RAND_1572 = {1{`RANDOM}};
  mesh_6_0_io_in_control_0_shift_pipe_b = _RAND_1572[4:0];
  _RAND_1573 = {1{`RANDOM}};
  mesh_6_0_io_in_control_0_dataflow_pipe_b = _RAND_1573[0:0];
  _RAND_1574 = {1{`RANDOM}};
  mesh_6_0_io_in_control_0_propagate_pipe_b = _RAND_1574[0:0];
  _RAND_1575 = {1{`RANDOM}};
  mesh_6_0_io_in_control_1_shift_pipe_b = _RAND_1575[4:0];
  _RAND_1576 = {1{`RANDOM}};
  mesh_6_0_io_in_control_1_dataflow_pipe_b = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  mesh_6_0_io_in_control_1_propagate_pipe_b = _RAND_1577[0:0];
  _RAND_1578 = {1{`RANDOM}};
  mesh_7_0_io_in_control_0_shift_pipe_b = _RAND_1578[4:0];
  _RAND_1579 = {1{`RANDOM}};
  mesh_7_0_io_in_control_0_dataflow_pipe_b = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  mesh_7_0_io_in_control_0_propagate_pipe_b = _RAND_1580[0:0];
  _RAND_1581 = {1{`RANDOM}};
  mesh_7_0_io_in_control_1_shift_pipe_b = _RAND_1581[4:0];
  _RAND_1582 = {1{`RANDOM}};
  mesh_7_0_io_in_control_1_dataflow_pipe_b = _RAND_1582[0:0];
  _RAND_1583 = {1{`RANDOM}};
  mesh_7_0_io_in_control_1_propagate_pipe_b = _RAND_1583[0:0];
  _RAND_1584 = {1{`RANDOM}};
  mesh_8_0_io_in_control_0_shift_pipe_b = _RAND_1584[4:0];
  _RAND_1585 = {1{`RANDOM}};
  mesh_8_0_io_in_control_0_dataflow_pipe_b = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  mesh_8_0_io_in_control_0_propagate_pipe_b = _RAND_1586[0:0];
  _RAND_1587 = {1{`RANDOM}};
  mesh_8_0_io_in_control_1_shift_pipe_b = _RAND_1587[4:0];
  _RAND_1588 = {1{`RANDOM}};
  mesh_8_0_io_in_control_1_dataflow_pipe_b = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  mesh_8_0_io_in_control_1_propagate_pipe_b = _RAND_1589[0:0];
  _RAND_1590 = {1{`RANDOM}};
  mesh_9_0_io_in_control_0_shift_pipe_b = _RAND_1590[4:0];
  _RAND_1591 = {1{`RANDOM}};
  mesh_9_0_io_in_control_0_dataflow_pipe_b = _RAND_1591[0:0];
  _RAND_1592 = {1{`RANDOM}};
  mesh_9_0_io_in_control_0_propagate_pipe_b = _RAND_1592[0:0];
  _RAND_1593 = {1{`RANDOM}};
  mesh_9_0_io_in_control_1_shift_pipe_b = _RAND_1593[4:0];
  _RAND_1594 = {1{`RANDOM}};
  mesh_9_0_io_in_control_1_dataflow_pipe_b = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  mesh_9_0_io_in_control_1_propagate_pipe_b = _RAND_1595[0:0];
  _RAND_1596 = {1{`RANDOM}};
  mesh_10_0_io_in_control_0_shift_pipe_b = _RAND_1596[4:0];
  _RAND_1597 = {1{`RANDOM}};
  mesh_10_0_io_in_control_0_dataflow_pipe_b = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  mesh_10_0_io_in_control_0_propagate_pipe_b = _RAND_1598[0:0];
  _RAND_1599 = {1{`RANDOM}};
  mesh_10_0_io_in_control_1_shift_pipe_b = _RAND_1599[4:0];
  _RAND_1600 = {1{`RANDOM}};
  mesh_10_0_io_in_control_1_dataflow_pipe_b = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  mesh_10_0_io_in_control_1_propagate_pipe_b = _RAND_1601[0:0];
  _RAND_1602 = {1{`RANDOM}};
  mesh_11_0_io_in_control_0_shift_pipe_b = _RAND_1602[4:0];
  _RAND_1603 = {1{`RANDOM}};
  mesh_11_0_io_in_control_0_dataflow_pipe_b = _RAND_1603[0:0];
  _RAND_1604 = {1{`RANDOM}};
  mesh_11_0_io_in_control_0_propagate_pipe_b = _RAND_1604[0:0];
  _RAND_1605 = {1{`RANDOM}};
  mesh_11_0_io_in_control_1_shift_pipe_b = _RAND_1605[4:0];
  _RAND_1606 = {1{`RANDOM}};
  mesh_11_0_io_in_control_1_dataflow_pipe_b = _RAND_1606[0:0];
  _RAND_1607 = {1{`RANDOM}};
  mesh_11_0_io_in_control_1_propagate_pipe_b = _RAND_1607[0:0];
  _RAND_1608 = {1{`RANDOM}};
  mesh_12_0_io_in_control_0_shift_pipe_b = _RAND_1608[4:0];
  _RAND_1609 = {1{`RANDOM}};
  mesh_12_0_io_in_control_0_dataflow_pipe_b = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  mesh_12_0_io_in_control_0_propagate_pipe_b = _RAND_1610[0:0];
  _RAND_1611 = {1{`RANDOM}};
  mesh_12_0_io_in_control_1_shift_pipe_b = _RAND_1611[4:0];
  _RAND_1612 = {1{`RANDOM}};
  mesh_12_0_io_in_control_1_dataflow_pipe_b = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  mesh_12_0_io_in_control_1_propagate_pipe_b = _RAND_1613[0:0];
  _RAND_1614 = {1{`RANDOM}};
  mesh_13_0_io_in_control_0_shift_pipe_b = _RAND_1614[4:0];
  _RAND_1615 = {1{`RANDOM}};
  mesh_13_0_io_in_control_0_dataflow_pipe_b = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  mesh_13_0_io_in_control_0_propagate_pipe_b = _RAND_1616[0:0];
  _RAND_1617 = {1{`RANDOM}};
  mesh_13_0_io_in_control_1_shift_pipe_b = _RAND_1617[4:0];
  _RAND_1618 = {1{`RANDOM}};
  mesh_13_0_io_in_control_1_dataflow_pipe_b = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  mesh_13_0_io_in_control_1_propagate_pipe_b = _RAND_1619[0:0];
  _RAND_1620 = {1{`RANDOM}};
  mesh_14_0_io_in_control_0_shift_pipe_b = _RAND_1620[4:0];
  _RAND_1621 = {1{`RANDOM}};
  mesh_14_0_io_in_control_0_dataflow_pipe_b = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  mesh_14_0_io_in_control_0_propagate_pipe_b = _RAND_1622[0:0];
  _RAND_1623 = {1{`RANDOM}};
  mesh_14_0_io_in_control_1_shift_pipe_b = _RAND_1623[4:0];
  _RAND_1624 = {1{`RANDOM}};
  mesh_14_0_io_in_control_1_dataflow_pipe_b = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  mesh_14_0_io_in_control_1_propagate_pipe_b = _RAND_1625[0:0];
  _RAND_1626 = {1{`RANDOM}};
  mesh_15_0_io_in_control_0_shift_pipe_b = _RAND_1626[4:0];
  _RAND_1627 = {1{`RANDOM}};
  mesh_15_0_io_in_control_0_dataflow_pipe_b = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  mesh_15_0_io_in_control_0_propagate_pipe_b = _RAND_1628[0:0];
  _RAND_1629 = {1{`RANDOM}};
  mesh_15_0_io_in_control_1_shift_pipe_b = _RAND_1629[4:0];
  _RAND_1630 = {1{`RANDOM}};
  mesh_15_0_io_in_control_1_dataflow_pipe_b = _RAND_1630[0:0];
  _RAND_1631 = {1{`RANDOM}};
  mesh_15_0_io_in_control_1_propagate_pipe_b = _RAND_1631[0:0];
  _RAND_1632 = {1{`RANDOM}};
  mesh_0_1_io_in_control_0_shift_pipe_b = _RAND_1632[4:0];
  _RAND_1633 = {1{`RANDOM}};
  mesh_0_1_io_in_control_0_dataflow_pipe_b = _RAND_1633[0:0];
  _RAND_1634 = {1{`RANDOM}};
  mesh_0_1_io_in_control_0_propagate_pipe_b = _RAND_1634[0:0];
  _RAND_1635 = {1{`RANDOM}};
  mesh_0_1_io_in_control_1_shift_pipe_b = _RAND_1635[4:0];
  _RAND_1636 = {1{`RANDOM}};
  mesh_0_1_io_in_control_1_dataflow_pipe_b = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  mesh_0_1_io_in_control_1_propagate_pipe_b = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  mesh_1_1_io_in_control_0_shift_pipe_b = _RAND_1638[4:0];
  _RAND_1639 = {1{`RANDOM}};
  mesh_1_1_io_in_control_0_dataflow_pipe_b = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  mesh_1_1_io_in_control_0_propagate_pipe_b = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  mesh_1_1_io_in_control_1_shift_pipe_b = _RAND_1641[4:0];
  _RAND_1642 = {1{`RANDOM}};
  mesh_1_1_io_in_control_1_dataflow_pipe_b = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  mesh_1_1_io_in_control_1_propagate_pipe_b = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  mesh_2_1_io_in_control_0_shift_pipe_b = _RAND_1644[4:0];
  _RAND_1645 = {1{`RANDOM}};
  mesh_2_1_io_in_control_0_dataflow_pipe_b = _RAND_1645[0:0];
  _RAND_1646 = {1{`RANDOM}};
  mesh_2_1_io_in_control_0_propagate_pipe_b = _RAND_1646[0:0];
  _RAND_1647 = {1{`RANDOM}};
  mesh_2_1_io_in_control_1_shift_pipe_b = _RAND_1647[4:0];
  _RAND_1648 = {1{`RANDOM}};
  mesh_2_1_io_in_control_1_dataflow_pipe_b = _RAND_1648[0:0];
  _RAND_1649 = {1{`RANDOM}};
  mesh_2_1_io_in_control_1_propagate_pipe_b = _RAND_1649[0:0];
  _RAND_1650 = {1{`RANDOM}};
  mesh_3_1_io_in_control_0_shift_pipe_b = _RAND_1650[4:0];
  _RAND_1651 = {1{`RANDOM}};
  mesh_3_1_io_in_control_0_dataflow_pipe_b = _RAND_1651[0:0];
  _RAND_1652 = {1{`RANDOM}};
  mesh_3_1_io_in_control_0_propagate_pipe_b = _RAND_1652[0:0];
  _RAND_1653 = {1{`RANDOM}};
  mesh_3_1_io_in_control_1_shift_pipe_b = _RAND_1653[4:0];
  _RAND_1654 = {1{`RANDOM}};
  mesh_3_1_io_in_control_1_dataflow_pipe_b = _RAND_1654[0:0];
  _RAND_1655 = {1{`RANDOM}};
  mesh_3_1_io_in_control_1_propagate_pipe_b = _RAND_1655[0:0];
  _RAND_1656 = {1{`RANDOM}};
  mesh_4_1_io_in_control_0_shift_pipe_b = _RAND_1656[4:0];
  _RAND_1657 = {1{`RANDOM}};
  mesh_4_1_io_in_control_0_dataflow_pipe_b = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  mesh_4_1_io_in_control_0_propagate_pipe_b = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  mesh_4_1_io_in_control_1_shift_pipe_b = _RAND_1659[4:0];
  _RAND_1660 = {1{`RANDOM}};
  mesh_4_1_io_in_control_1_dataflow_pipe_b = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  mesh_4_1_io_in_control_1_propagate_pipe_b = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  mesh_5_1_io_in_control_0_shift_pipe_b = _RAND_1662[4:0];
  _RAND_1663 = {1{`RANDOM}};
  mesh_5_1_io_in_control_0_dataflow_pipe_b = _RAND_1663[0:0];
  _RAND_1664 = {1{`RANDOM}};
  mesh_5_1_io_in_control_0_propagate_pipe_b = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  mesh_5_1_io_in_control_1_shift_pipe_b = _RAND_1665[4:0];
  _RAND_1666 = {1{`RANDOM}};
  mesh_5_1_io_in_control_1_dataflow_pipe_b = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  mesh_5_1_io_in_control_1_propagate_pipe_b = _RAND_1667[0:0];
  _RAND_1668 = {1{`RANDOM}};
  mesh_6_1_io_in_control_0_shift_pipe_b = _RAND_1668[4:0];
  _RAND_1669 = {1{`RANDOM}};
  mesh_6_1_io_in_control_0_dataflow_pipe_b = _RAND_1669[0:0];
  _RAND_1670 = {1{`RANDOM}};
  mesh_6_1_io_in_control_0_propagate_pipe_b = _RAND_1670[0:0];
  _RAND_1671 = {1{`RANDOM}};
  mesh_6_1_io_in_control_1_shift_pipe_b = _RAND_1671[4:0];
  _RAND_1672 = {1{`RANDOM}};
  mesh_6_1_io_in_control_1_dataflow_pipe_b = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  mesh_6_1_io_in_control_1_propagate_pipe_b = _RAND_1673[0:0];
  _RAND_1674 = {1{`RANDOM}};
  mesh_7_1_io_in_control_0_shift_pipe_b = _RAND_1674[4:0];
  _RAND_1675 = {1{`RANDOM}};
  mesh_7_1_io_in_control_0_dataflow_pipe_b = _RAND_1675[0:0];
  _RAND_1676 = {1{`RANDOM}};
  mesh_7_1_io_in_control_0_propagate_pipe_b = _RAND_1676[0:0];
  _RAND_1677 = {1{`RANDOM}};
  mesh_7_1_io_in_control_1_shift_pipe_b = _RAND_1677[4:0];
  _RAND_1678 = {1{`RANDOM}};
  mesh_7_1_io_in_control_1_dataflow_pipe_b = _RAND_1678[0:0];
  _RAND_1679 = {1{`RANDOM}};
  mesh_7_1_io_in_control_1_propagate_pipe_b = _RAND_1679[0:0];
  _RAND_1680 = {1{`RANDOM}};
  mesh_8_1_io_in_control_0_shift_pipe_b = _RAND_1680[4:0];
  _RAND_1681 = {1{`RANDOM}};
  mesh_8_1_io_in_control_0_dataflow_pipe_b = _RAND_1681[0:0];
  _RAND_1682 = {1{`RANDOM}};
  mesh_8_1_io_in_control_0_propagate_pipe_b = _RAND_1682[0:0];
  _RAND_1683 = {1{`RANDOM}};
  mesh_8_1_io_in_control_1_shift_pipe_b = _RAND_1683[4:0];
  _RAND_1684 = {1{`RANDOM}};
  mesh_8_1_io_in_control_1_dataflow_pipe_b = _RAND_1684[0:0];
  _RAND_1685 = {1{`RANDOM}};
  mesh_8_1_io_in_control_1_propagate_pipe_b = _RAND_1685[0:0];
  _RAND_1686 = {1{`RANDOM}};
  mesh_9_1_io_in_control_0_shift_pipe_b = _RAND_1686[4:0];
  _RAND_1687 = {1{`RANDOM}};
  mesh_9_1_io_in_control_0_dataflow_pipe_b = _RAND_1687[0:0];
  _RAND_1688 = {1{`RANDOM}};
  mesh_9_1_io_in_control_0_propagate_pipe_b = _RAND_1688[0:0];
  _RAND_1689 = {1{`RANDOM}};
  mesh_9_1_io_in_control_1_shift_pipe_b = _RAND_1689[4:0];
  _RAND_1690 = {1{`RANDOM}};
  mesh_9_1_io_in_control_1_dataflow_pipe_b = _RAND_1690[0:0];
  _RAND_1691 = {1{`RANDOM}};
  mesh_9_1_io_in_control_1_propagate_pipe_b = _RAND_1691[0:0];
  _RAND_1692 = {1{`RANDOM}};
  mesh_10_1_io_in_control_0_shift_pipe_b = _RAND_1692[4:0];
  _RAND_1693 = {1{`RANDOM}};
  mesh_10_1_io_in_control_0_dataflow_pipe_b = _RAND_1693[0:0];
  _RAND_1694 = {1{`RANDOM}};
  mesh_10_1_io_in_control_0_propagate_pipe_b = _RAND_1694[0:0];
  _RAND_1695 = {1{`RANDOM}};
  mesh_10_1_io_in_control_1_shift_pipe_b = _RAND_1695[4:0];
  _RAND_1696 = {1{`RANDOM}};
  mesh_10_1_io_in_control_1_dataflow_pipe_b = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  mesh_10_1_io_in_control_1_propagate_pipe_b = _RAND_1697[0:0];
  _RAND_1698 = {1{`RANDOM}};
  mesh_11_1_io_in_control_0_shift_pipe_b = _RAND_1698[4:0];
  _RAND_1699 = {1{`RANDOM}};
  mesh_11_1_io_in_control_0_dataflow_pipe_b = _RAND_1699[0:0];
  _RAND_1700 = {1{`RANDOM}};
  mesh_11_1_io_in_control_0_propagate_pipe_b = _RAND_1700[0:0];
  _RAND_1701 = {1{`RANDOM}};
  mesh_11_1_io_in_control_1_shift_pipe_b = _RAND_1701[4:0];
  _RAND_1702 = {1{`RANDOM}};
  mesh_11_1_io_in_control_1_dataflow_pipe_b = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  mesh_11_1_io_in_control_1_propagate_pipe_b = _RAND_1703[0:0];
  _RAND_1704 = {1{`RANDOM}};
  mesh_12_1_io_in_control_0_shift_pipe_b = _RAND_1704[4:0];
  _RAND_1705 = {1{`RANDOM}};
  mesh_12_1_io_in_control_0_dataflow_pipe_b = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  mesh_12_1_io_in_control_0_propagate_pipe_b = _RAND_1706[0:0];
  _RAND_1707 = {1{`RANDOM}};
  mesh_12_1_io_in_control_1_shift_pipe_b = _RAND_1707[4:0];
  _RAND_1708 = {1{`RANDOM}};
  mesh_12_1_io_in_control_1_dataflow_pipe_b = _RAND_1708[0:0];
  _RAND_1709 = {1{`RANDOM}};
  mesh_12_1_io_in_control_1_propagate_pipe_b = _RAND_1709[0:0];
  _RAND_1710 = {1{`RANDOM}};
  mesh_13_1_io_in_control_0_shift_pipe_b = _RAND_1710[4:0];
  _RAND_1711 = {1{`RANDOM}};
  mesh_13_1_io_in_control_0_dataflow_pipe_b = _RAND_1711[0:0];
  _RAND_1712 = {1{`RANDOM}};
  mesh_13_1_io_in_control_0_propagate_pipe_b = _RAND_1712[0:0];
  _RAND_1713 = {1{`RANDOM}};
  mesh_13_1_io_in_control_1_shift_pipe_b = _RAND_1713[4:0];
  _RAND_1714 = {1{`RANDOM}};
  mesh_13_1_io_in_control_1_dataflow_pipe_b = _RAND_1714[0:0];
  _RAND_1715 = {1{`RANDOM}};
  mesh_13_1_io_in_control_1_propagate_pipe_b = _RAND_1715[0:0];
  _RAND_1716 = {1{`RANDOM}};
  mesh_14_1_io_in_control_0_shift_pipe_b = _RAND_1716[4:0];
  _RAND_1717 = {1{`RANDOM}};
  mesh_14_1_io_in_control_0_dataflow_pipe_b = _RAND_1717[0:0];
  _RAND_1718 = {1{`RANDOM}};
  mesh_14_1_io_in_control_0_propagate_pipe_b = _RAND_1718[0:0];
  _RAND_1719 = {1{`RANDOM}};
  mesh_14_1_io_in_control_1_shift_pipe_b = _RAND_1719[4:0];
  _RAND_1720 = {1{`RANDOM}};
  mesh_14_1_io_in_control_1_dataflow_pipe_b = _RAND_1720[0:0];
  _RAND_1721 = {1{`RANDOM}};
  mesh_14_1_io_in_control_1_propagate_pipe_b = _RAND_1721[0:0];
  _RAND_1722 = {1{`RANDOM}};
  mesh_15_1_io_in_control_0_shift_pipe_b = _RAND_1722[4:0];
  _RAND_1723 = {1{`RANDOM}};
  mesh_15_1_io_in_control_0_dataflow_pipe_b = _RAND_1723[0:0];
  _RAND_1724 = {1{`RANDOM}};
  mesh_15_1_io_in_control_0_propagate_pipe_b = _RAND_1724[0:0];
  _RAND_1725 = {1{`RANDOM}};
  mesh_15_1_io_in_control_1_shift_pipe_b = _RAND_1725[4:0];
  _RAND_1726 = {1{`RANDOM}};
  mesh_15_1_io_in_control_1_dataflow_pipe_b = _RAND_1726[0:0];
  _RAND_1727 = {1{`RANDOM}};
  mesh_15_1_io_in_control_1_propagate_pipe_b = _RAND_1727[0:0];
  _RAND_1728 = {1{`RANDOM}};
  mesh_0_2_io_in_control_0_shift_pipe_b = _RAND_1728[4:0];
  _RAND_1729 = {1{`RANDOM}};
  mesh_0_2_io_in_control_0_dataflow_pipe_b = _RAND_1729[0:0];
  _RAND_1730 = {1{`RANDOM}};
  mesh_0_2_io_in_control_0_propagate_pipe_b = _RAND_1730[0:0];
  _RAND_1731 = {1{`RANDOM}};
  mesh_0_2_io_in_control_1_shift_pipe_b = _RAND_1731[4:0];
  _RAND_1732 = {1{`RANDOM}};
  mesh_0_2_io_in_control_1_dataflow_pipe_b = _RAND_1732[0:0];
  _RAND_1733 = {1{`RANDOM}};
  mesh_0_2_io_in_control_1_propagate_pipe_b = _RAND_1733[0:0];
  _RAND_1734 = {1{`RANDOM}};
  mesh_1_2_io_in_control_0_shift_pipe_b = _RAND_1734[4:0];
  _RAND_1735 = {1{`RANDOM}};
  mesh_1_2_io_in_control_0_dataflow_pipe_b = _RAND_1735[0:0];
  _RAND_1736 = {1{`RANDOM}};
  mesh_1_2_io_in_control_0_propagate_pipe_b = _RAND_1736[0:0];
  _RAND_1737 = {1{`RANDOM}};
  mesh_1_2_io_in_control_1_shift_pipe_b = _RAND_1737[4:0];
  _RAND_1738 = {1{`RANDOM}};
  mesh_1_2_io_in_control_1_dataflow_pipe_b = _RAND_1738[0:0];
  _RAND_1739 = {1{`RANDOM}};
  mesh_1_2_io_in_control_1_propagate_pipe_b = _RAND_1739[0:0];
  _RAND_1740 = {1{`RANDOM}};
  mesh_2_2_io_in_control_0_shift_pipe_b = _RAND_1740[4:0];
  _RAND_1741 = {1{`RANDOM}};
  mesh_2_2_io_in_control_0_dataflow_pipe_b = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  mesh_2_2_io_in_control_0_propagate_pipe_b = _RAND_1742[0:0];
  _RAND_1743 = {1{`RANDOM}};
  mesh_2_2_io_in_control_1_shift_pipe_b = _RAND_1743[4:0];
  _RAND_1744 = {1{`RANDOM}};
  mesh_2_2_io_in_control_1_dataflow_pipe_b = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  mesh_2_2_io_in_control_1_propagate_pipe_b = _RAND_1745[0:0];
  _RAND_1746 = {1{`RANDOM}};
  mesh_3_2_io_in_control_0_shift_pipe_b = _RAND_1746[4:0];
  _RAND_1747 = {1{`RANDOM}};
  mesh_3_2_io_in_control_0_dataflow_pipe_b = _RAND_1747[0:0];
  _RAND_1748 = {1{`RANDOM}};
  mesh_3_2_io_in_control_0_propagate_pipe_b = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  mesh_3_2_io_in_control_1_shift_pipe_b = _RAND_1749[4:0];
  _RAND_1750 = {1{`RANDOM}};
  mesh_3_2_io_in_control_1_dataflow_pipe_b = _RAND_1750[0:0];
  _RAND_1751 = {1{`RANDOM}};
  mesh_3_2_io_in_control_1_propagate_pipe_b = _RAND_1751[0:0];
  _RAND_1752 = {1{`RANDOM}};
  mesh_4_2_io_in_control_0_shift_pipe_b = _RAND_1752[4:0];
  _RAND_1753 = {1{`RANDOM}};
  mesh_4_2_io_in_control_0_dataflow_pipe_b = _RAND_1753[0:0];
  _RAND_1754 = {1{`RANDOM}};
  mesh_4_2_io_in_control_0_propagate_pipe_b = _RAND_1754[0:0];
  _RAND_1755 = {1{`RANDOM}};
  mesh_4_2_io_in_control_1_shift_pipe_b = _RAND_1755[4:0];
  _RAND_1756 = {1{`RANDOM}};
  mesh_4_2_io_in_control_1_dataflow_pipe_b = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  mesh_4_2_io_in_control_1_propagate_pipe_b = _RAND_1757[0:0];
  _RAND_1758 = {1{`RANDOM}};
  mesh_5_2_io_in_control_0_shift_pipe_b = _RAND_1758[4:0];
  _RAND_1759 = {1{`RANDOM}};
  mesh_5_2_io_in_control_0_dataflow_pipe_b = _RAND_1759[0:0];
  _RAND_1760 = {1{`RANDOM}};
  mesh_5_2_io_in_control_0_propagate_pipe_b = _RAND_1760[0:0];
  _RAND_1761 = {1{`RANDOM}};
  mesh_5_2_io_in_control_1_shift_pipe_b = _RAND_1761[4:0];
  _RAND_1762 = {1{`RANDOM}};
  mesh_5_2_io_in_control_1_dataflow_pipe_b = _RAND_1762[0:0];
  _RAND_1763 = {1{`RANDOM}};
  mesh_5_2_io_in_control_1_propagate_pipe_b = _RAND_1763[0:0];
  _RAND_1764 = {1{`RANDOM}};
  mesh_6_2_io_in_control_0_shift_pipe_b = _RAND_1764[4:0];
  _RAND_1765 = {1{`RANDOM}};
  mesh_6_2_io_in_control_0_dataflow_pipe_b = _RAND_1765[0:0];
  _RAND_1766 = {1{`RANDOM}};
  mesh_6_2_io_in_control_0_propagate_pipe_b = _RAND_1766[0:0];
  _RAND_1767 = {1{`RANDOM}};
  mesh_6_2_io_in_control_1_shift_pipe_b = _RAND_1767[4:0];
  _RAND_1768 = {1{`RANDOM}};
  mesh_6_2_io_in_control_1_dataflow_pipe_b = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  mesh_6_2_io_in_control_1_propagate_pipe_b = _RAND_1769[0:0];
  _RAND_1770 = {1{`RANDOM}};
  mesh_7_2_io_in_control_0_shift_pipe_b = _RAND_1770[4:0];
  _RAND_1771 = {1{`RANDOM}};
  mesh_7_2_io_in_control_0_dataflow_pipe_b = _RAND_1771[0:0];
  _RAND_1772 = {1{`RANDOM}};
  mesh_7_2_io_in_control_0_propagate_pipe_b = _RAND_1772[0:0];
  _RAND_1773 = {1{`RANDOM}};
  mesh_7_2_io_in_control_1_shift_pipe_b = _RAND_1773[4:0];
  _RAND_1774 = {1{`RANDOM}};
  mesh_7_2_io_in_control_1_dataflow_pipe_b = _RAND_1774[0:0];
  _RAND_1775 = {1{`RANDOM}};
  mesh_7_2_io_in_control_1_propagate_pipe_b = _RAND_1775[0:0];
  _RAND_1776 = {1{`RANDOM}};
  mesh_8_2_io_in_control_0_shift_pipe_b = _RAND_1776[4:0];
  _RAND_1777 = {1{`RANDOM}};
  mesh_8_2_io_in_control_0_dataflow_pipe_b = _RAND_1777[0:0];
  _RAND_1778 = {1{`RANDOM}};
  mesh_8_2_io_in_control_0_propagate_pipe_b = _RAND_1778[0:0];
  _RAND_1779 = {1{`RANDOM}};
  mesh_8_2_io_in_control_1_shift_pipe_b = _RAND_1779[4:0];
  _RAND_1780 = {1{`RANDOM}};
  mesh_8_2_io_in_control_1_dataflow_pipe_b = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  mesh_8_2_io_in_control_1_propagate_pipe_b = _RAND_1781[0:0];
  _RAND_1782 = {1{`RANDOM}};
  mesh_9_2_io_in_control_0_shift_pipe_b = _RAND_1782[4:0];
  _RAND_1783 = {1{`RANDOM}};
  mesh_9_2_io_in_control_0_dataflow_pipe_b = _RAND_1783[0:0];
  _RAND_1784 = {1{`RANDOM}};
  mesh_9_2_io_in_control_0_propagate_pipe_b = _RAND_1784[0:0];
  _RAND_1785 = {1{`RANDOM}};
  mesh_9_2_io_in_control_1_shift_pipe_b = _RAND_1785[4:0];
  _RAND_1786 = {1{`RANDOM}};
  mesh_9_2_io_in_control_1_dataflow_pipe_b = _RAND_1786[0:0];
  _RAND_1787 = {1{`RANDOM}};
  mesh_9_2_io_in_control_1_propagate_pipe_b = _RAND_1787[0:0];
  _RAND_1788 = {1{`RANDOM}};
  mesh_10_2_io_in_control_0_shift_pipe_b = _RAND_1788[4:0];
  _RAND_1789 = {1{`RANDOM}};
  mesh_10_2_io_in_control_0_dataflow_pipe_b = _RAND_1789[0:0];
  _RAND_1790 = {1{`RANDOM}};
  mesh_10_2_io_in_control_0_propagate_pipe_b = _RAND_1790[0:0];
  _RAND_1791 = {1{`RANDOM}};
  mesh_10_2_io_in_control_1_shift_pipe_b = _RAND_1791[4:0];
  _RAND_1792 = {1{`RANDOM}};
  mesh_10_2_io_in_control_1_dataflow_pipe_b = _RAND_1792[0:0];
  _RAND_1793 = {1{`RANDOM}};
  mesh_10_2_io_in_control_1_propagate_pipe_b = _RAND_1793[0:0];
  _RAND_1794 = {1{`RANDOM}};
  mesh_11_2_io_in_control_0_shift_pipe_b = _RAND_1794[4:0];
  _RAND_1795 = {1{`RANDOM}};
  mesh_11_2_io_in_control_0_dataflow_pipe_b = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  mesh_11_2_io_in_control_0_propagate_pipe_b = _RAND_1796[0:0];
  _RAND_1797 = {1{`RANDOM}};
  mesh_11_2_io_in_control_1_shift_pipe_b = _RAND_1797[4:0];
  _RAND_1798 = {1{`RANDOM}};
  mesh_11_2_io_in_control_1_dataflow_pipe_b = _RAND_1798[0:0];
  _RAND_1799 = {1{`RANDOM}};
  mesh_11_2_io_in_control_1_propagate_pipe_b = _RAND_1799[0:0];
  _RAND_1800 = {1{`RANDOM}};
  mesh_12_2_io_in_control_0_shift_pipe_b = _RAND_1800[4:0];
  _RAND_1801 = {1{`RANDOM}};
  mesh_12_2_io_in_control_0_dataflow_pipe_b = _RAND_1801[0:0];
  _RAND_1802 = {1{`RANDOM}};
  mesh_12_2_io_in_control_0_propagate_pipe_b = _RAND_1802[0:0];
  _RAND_1803 = {1{`RANDOM}};
  mesh_12_2_io_in_control_1_shift_pipe_b = _RAND_1803[4:0];
  _RAND_1804 = {1{`RANDOM}};
  mesh_12_2_io_in_control_1_dataflow_pipe_b = _RAND_1804[0:0];
  _RAND_1805 = {1{`RANDOM}};
  mesh_12_2_io_in_control_1_propagate_pipe_b = _RAND_1805[0:0];
  _RAND_1806 = {1{`RANDOM}};
  mesh_13_2_io_in_control_0_shift_pipe_b = _RAND_1806[4:0];
  _RAND_1807 = {1{`RANDOM}};
  mesh_13_2_io_in_control_0_dataflow_pipe_b = _RAND_1807[0:0];
  _RAND_1808 = {1{`RANDOM}};
  mesh_13_2_io_in_control_0_propagate_pipe_b = _RAND_1808[0:0];
  _RAND_1809 = {1{`RANDOM}};
  mesh_13_2_io_in_control_1_shift_pipe_b = _RAND_1809[4:0];
  _RAND_1810 = {1{`RANDOM}};
  mesh_13_2_io_in_control_1_dataflow_pipe_b = _RAND_1810[0:0];
  _RAND_1811 = {1{`RANDOM}};
  mesh_13_2_io_in_control_1_propagate_pipe_b = _RAND_1811[0:0];
  _RAND_1812 = {1{`RANDOM}};
  mesh_14_2_io_in_control_0_shift_pipe_b = _RAND_1812[4:0];
  _RAND_1813 = {1{`RANDOM}};
  mesh_14_2_io_in_control_0_dataflow_pipe_b = _RAND_1813[0:0];
  _RAND_1814 = {1{`RANDOM}};
  mesh_14_2_io_in_control_0_propagate_pipe_b = _RAND_1814[0:0];
  _RAND_1815 = {1{`RANDOM}};
  mesh_14_2_io_in_control_1_shift_pipe_b = _RAND_1815[4:0];
  _RAND_1816 = {1{`RANDOM}};
  mesh_14_2_io_in_control_1_dataflow_pipe_b = _RAND_1816[0:0];
  _RAND_1817 = {1{`RANDOM}};
  mesh_14_2_io_in_control_1_propagate_pipe_b = _RAND_1817[0:0];
  _RAND_1818 = {1{`RANDOM}};
  mesh_15_2_io_in_control_0_shift_pipe_b = _RAND_1818[4:0];
  _RAND_1819 = {1{`RANDOM}};
  mesh_15_2_io_in_control_0_dataflow_pipe_b = _RAND_1819[0:0];
  _RAND_1820 = {1{`RANDOM}};
  mesh_15_2_io_in_control_0_propagate_pipe_b = _RAND_1820[0:0];
  _RAND_1821 = {1{`RANDOM}};
  mesh_15_2_io_in_control_1_shift_pipe_b = _RAND_1821[4:0];
  _RAND_1822 = {1{`RANDOM}};
  mesh_15_2_io_in_control_1_dataflow_pipe_b = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  mesh_15_2_io_in_control_1_propagate_pipe_b = _RAND_1823[0:0];
  _RAND_1824 = {1{`RANDOM}};
  mesh_0_3_io_in_control_0_shift_pipe_b = _RAND_1824[4:0];
  _RAND_1825 = {1{`RANDOM}};
  mesh_0_3_io_in_control_0_dataflow_pipe_b = _RAND_1825[0:0];
  _RAND_1826 = {1{`RANDOM}};
  mesh_0_3_io_in_control_0_propagate_pipe_b = _RAND_1826[0:0];
  _RAND_1827 = {1{`RANDOM}};
  mesh_0_3_io_in_control_1_shift_pipe_b = _RAND_1827[4:0];
  _RAND_1828 = {1{`RANDOM}};
  mesh_0_3_io_in_control_1_dataflow_pipe_b = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  mesh_0_3_io_in_control_1_propagate_pipe_b = _RAND_1829[0:0];
  _RAND_1830 = {1{`RANDOM}};
  mesh_1_3_io_in_control_0_shift_pipe_b = _RAND_1830[4:0];
  _RAND_1831 = {1{`RANDOM}};
  mesh_1_3_io_in_control_0_dataflow_pipe_b = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  mesh_1_3_io_in_control_0_propagate_pipe_b = _RAND_1832[0:0];
  _RAND_1833 = {1{`RANDOM}};
  mesh_1_3_io_in_control_1_shift_pipe_b = _RAND_1833[4:0];
  _RAND_1834 = {1{`RANDOM}};
  mesh_1_3_io_in_control_1_dataflow_pipe_b = _RAND_1834[0:0];
  _RAND_1835 = {1{`RANDOM}};
  mesh_1_3_io_in_control_1_propagate_pipe_b = _RAND_1835[0:0];
  _RAND_1836 = {1{`RANDOM}};
  mesh_2_3_io_in_control_0_shift_pipe_b = _RAND_1836[4:0];
  _RAND_1837 = {1{`RANDOM}};
  mesh_2_3_io_in_control_0_dataflow_pipe_b = _RAND_1837[0:0];
  _RAND_1838 = {1{`RANDOM}};
  mesh_2_3_io_in_control_0_propagate_pipe_b = _RAND_1838[0:0];
  _RAND_1839 = {1{`RANDOM}};
  mesh_2_3_io_in_control_1_shift_pipe_b = _RAND_1839[4:0];
  _RAND_1840 = {1{`RANDOM}};
  mesh_2_3_io_in_control_1_dataflow_pipe_b = _RAND_1840[0:0];
  _RAND_1841 = {1{`RANDOM}};
  mesh_2_3_io_in_control_1_propagate_pipe_b = _RAND_1841[0:0];
  _RAND_1842 = {1{`RANDOM}};
  mesh_3_3_io_in_control_0_shift_pipe_b = _RAND_1842[4:0];
  _RAND_1843 = {1{`RANDOM}};
  mesh_3_3_io_in_control_0_dataflow_pipe_b = _RAND_1843[0:0];
  _RAND_1844 = {1{`RANDOM}};
  mesh_3_3_io_in_control_0_propagate_pipe_b = _RAND_1844[0:0];
  _RAND_1845 = {1{`RANDOM}};
  mesh_3_3_io_in_control_1_shift_pipe_b = _RAND_1845[4:0];
  _RAND_1846 = {1{`RANDOM}};
  mesh_3_3_io_in_control_1_dataflow_pipe_b = _RAND_1846[0:0];
  _RAND_1847 = {1{`RANDOM}};
  mesh_3_3_io_in_control_1_propagate_pipe_b = _RAND_1847[0:0];
  _RAND_1848 = {1{`RANDOM}};
  mesh_4_3_io_in_control_0_shift_pipe_b = _RAND_1848[4:0];
  _RAND_1849 = {1{`RANDOM}};
  mesh_4_3_io_in_control_0_dataflow_pipe_b = _RAND_1849[0:0];
  _RAND_1850 = {1{`RANDOM}};
  mesh_4_3_io_in_control_0_propagate_pipe_b = _RAND_1850[0:0];
  _RAND_1851 = {1{`RANDOM}};
  mesh_4_3_io_in_control_1_shift_pipe_b = _RAND_1851[4:0];
  _RAND_1852 = {1{`RANDOM}};
  mesh_4_3_io_in_control_1_dataflow_pipe_b = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  mesh_4_3_io_in_control_1_propagate_pipe_b = _RAND_1853[0:0];
  _RAND_1854 = {1{`RANDOM}};
  mesh_5_3_io_in_control_0_shift_pipe_b = _RAND_1854[4:0];
  _RAND_1855 = {1{`RANDOM}};
  mesh_5_3_io_in_control_0_dataflow_pipe_b = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  mesh_5_3_io_in_control_0_propagate_pipe_b = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  mesh_5_3_io_in_control_1_shift_pipe_b = _RAND_1857[4:0];
  _RAND_1858 = {1{`RANDOM}};
  mesh_5_3_io_in_control_1_dataflow_pipe_b = _RAND_1858[0:0];
  _RAND_1859 = {1{`RANDOM}};
  mesh_5_3_io_in_control_1_propagate_pipe_b = _RAND_1859[0:0];
  _RAND_1860 = {1{`RANDOM}};
  mesh_6_3_io_in_control_0_shift_pipe_b = _RAND_1860[4:0];
  _RAND_1861 = {1{`RANDOM}};
  mesh_6_3_io_in_control_0_dataflow_pipe_b = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  mesh_6_3_io_in_control_0_propagate_pipe_b = _RAND_1862[0:0];
  _RAND_1863 = {1{`RANDOM}};
  mesh_6_3_io_in_control_1_shift_pipe_b = _RAND_1863[4:0];
  _RAND_1864 = {1{`RANDOM}};
  mesh_6_3_io_in_control_1_dataflow_pipe_b = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  mesh_6_3_io_in_control_1_propagate_pipe_b = _RAND_1865[0:0];
  _RAND_1866 = {1{`RANDOM}};
  mesh_7_3_io_in_control_0_shift_pipe_b = _RAND_1866[4:0];
  _RAND_1867 = {1{`RANDOM}};
  mesh_7_3_io_in_control_0_dataflow_pipe_b = _RAND_1867[0:0];
  _RAND_1868 = {1{`RANDOM}};
  mesh_7_3_io_in_control_0_propagate_pipe_b = _RAND_1868[0:0];
  _RAND_1869 = {1{`RANDOM}};
  mesh_7_3_io_in_control_1_shift_pipe_b = _RAND_1869[4:0];
  _RAND_1870 = {1{`RANDOM}};
  mesh_7_3_io_in_control_1_dataflow_pipe_b = _RAND_1870[0:0];
  _RAND_1871 = {1{`RANDOM}};
  mesh_7_3_io_in_control_1_propagate_pipe_b = _RAND_1871[0:0];
  _RAND_1872 = {1{`RANDOM}};
  mesh_8_3_io_in_control_0_shift_pipe_b = _RAND_1872[4:0];
  _RAND_1873 = {1{`RANDOM}};
  mesh_8_3_io_in_control_0_dataflow_pipe_b = _RAND_1873[0:0];
  _RAND_1874 = {1{`RANDOM}};
  mesh_8_3_io_in_control_0_propagate_pipe_b = _RAND_1874[0:0];
  _RAND_1875 = {1{`RANDOM}};
  mesh_8_3_io_in_control_1_shift_pipe_b = _RAND_1875[4:0];
  _RAND_1876 = {1{`RANDOM}};
  mesh_8_3_io_in_control_1_dataflow_pipe_b = _RAND_1876[0:0];
  _RAND_1877 = {1{`RANDOM}};
  mesh_8_3_io_in_control_1_propagate_pipe_b = _RAND_1877[0:0];
  _RAND_1878 = {1{`RANDOM}};
  mesh_9_3_io_in_control_0_shift_pipe_b = _RAND_1878[4:0];
  _RAND_1879 = {1{`RANDOM}};
  mesh_9_3_io_in_control_0_dataflow_pipe_b = _RAND_1879[0:0];
  _RAND_1880 = {1{`RANDOM}};
  mesh_9_3_io_in_control_0_propagate_pipe_b = _RAND_1880[0:0];
  _RAND_1881 = {1{`RANDOM}};
  mesh_9_3_io_in_control_1_shift_pipe_b = _RAND_1881[4:0];
  _RAND_1882 = {1{`RANDOM}};
  mesh_9_3_io_in_control_1_dataflow_pipe_b = _RAND_1882[0:0];
  _RAND_1883 = {1{`RANDOM}};
  mesh_9_3_io_in_control_1_propagate_pipe_b = _RAND_1883[0:0];
  _RAND_1884 = {1{`RANDOM}};
  mesh_10_3_io_in_control_0_shift_pipe_b = _RAND_1884[4:0];
  _RAND_1885 = {1{`RANDOM}};
  mesh_10_3_io_in_control_0_dataflow_pipe_b = _RAND_1885[0:0];
  _RAND_1886 = {1{`RANDOM}};
  mesh_10_3_io_in_control_0_propagate_pipe_b = _RAND_1886[0:0];
  _RAND_1887 = {1{`RANDOM}};
  mesh_10_3_io_in_control_1_shift_pipe_b = _RAND_1887[4:0];
  _RAND_1888 = {1{`RANDOM}};
  mesh_10_3_io_in_control_1_dataflow_pipe_b = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  mesh_10_3_io_in_control_1_propagate_pipe_b = _RAND_1889[0:0];
  _RAND_1890 = {1{`RANDOM}};
  mesh_11_3_io_in_control_0_shift_pipe_b = _RAND_1890[4:0];
  _RAND_1891 = {1{`RANDOM}};
  mesh_11_3_io_in_control_0_dataflow_pipe_b = _RAND_1891[0:0];
  _RAND_1892 = {1{`RANDOM}};
  mesh_11_3_io_in_control_0_propagate_pipe_b = _RAND_1892[0:0];
  _RAND_1893 = {1{`RANDOM}};
  mesh_11_3_io_in_control_1_shift_pipe_b = _RAND_1893[4:0];
  _RAND_1894 = {1{`RANDOM}};
  mesh_11_3_io_in_control_1_dataflow_pipe_b = _RAND_1894[0:0];
  _RAND_1895 = {1{`RANDOM}};
  mesh_11_3_io_in_control_1_propagate_pipe_b = _RAND_1895[0:0];
  _RAND_1896 = {1{`RANDOM}};
  mesh_12_3_io_in_control_0_shift_pipe_b = _RAND_1896[4:0];
  _RAND_1897 = {1{`RANDOM}};
  mesh_12_3_io_in_control_0_dataflow_pipe_b = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  mesh_12_3_io_in_control_0_propagate_pipe_b = _RAND_1898[0:0];
  _RAND_1899 = {1{`RANDOM}};
  mesh_12_3_io_in_control_1_shift_pipe_b = _RAND_1899[4:0];
  _RAND_1900 = {1{`RANDOM}};
  mesh_12_3_io_in_control_1_dataflow_pipe_b = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  mesh_12_3_io_in_control_1_propagate_pipe_b = _RAND_1901[0:0];
  _RAND_1902 = {1{`RANDOM}};
  mesh_13_3_io_in_control_0_shift_pipe_b = _RAND_1902[4:0];
  _RAND_1903 = {1{`RANDOM}};
  mesh_13_3_io_in_control_0_dataflow_pipe_b = _RAND_1903[0:0];
  _RAND_1904 = {1{`RANDOM}};
  mesh_13_3_io_in_control_0_propagate_pipe_b = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  mesh_13_3_io_in_control_1_shift_pipe_b = _RAND_1905[4:0];
  _RAND_1906 = {1{`RANDOM}};
  mesh_13_3_io_in_control_1_dataflow_pipe_b = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  mesh_13_3_io_in_control_1_propagate_pipe_b = _RAND_1907[0:0];
  _RAND_1908 = {1{`RANDOM}};
  mesh_14_3_io_in_control_0_shift_pipe_b = _RAND_1908[4:0];
  _RAND_1909 = {1{`RANDOM}};
  mesh_14_3_io_in_control_0_dataflow_pipe_b = _RAND_1909[0:0];
  _RAND_1910 = {1{`RANDOM}};
  mesh_14_3_io_in_control_0_propagate_pipe_b = _RAND_1910[0:0];
  _RAND_1911 = {1{`RANDOM}};
  mesh_14_3_io_in_control_1_shift_pipe_b = _RAND_1911[4:0];
  _RAND_1912 = {1{`RANDOM}};
  mesh_14_3_io_in_control_1_dataflow_pipe_b = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  mesh_14_3_io_in_control_1_propagate_pipe_b = _RAND_1913[0:0];
  _RAND_1914 = {1{`RANDOM}};
  mesh_15_3_io_in_control_0_shift_pipe_b = _RAND_1914[4:0];
  _RAND_1915 = {1{`RANDOM}};
  mesh_15_3_io_in_control_0_dataflow_pipe_b = _RAND_1915[0:0];
  _RAND_1916 = {1{`RANDOM}};
  mesh_15_3_io_in_control_0_propagate_pipe_b = _RAND_1916[0:0];
  _RAND_1917 = {1{`RANDOM}};
  mesh_15_3_io_in_control_1_shift_pipe_b = _RAND_1917[4:0];
  _RAND_1918 = {1{`RANDOM}};
  mesh_15_3_io_in_control_1_dataflow_pipe_b = _RAND_1918[0:0];
  _RAND_1919 = {1{`RANDOM}};
  mesh_15_3_io_in_control_1_propagate_pipe_b = _RAND_1919[0:0];
  _RAND_1920 = {1{`RANDOM}};
  mesh_0_4_io_in_control_0_shift_pipe_b = _RAND_1920[4:0];
  _RAND_1921 = {1{`RANDOM}};
  mesh_0_4_io_in_control_0_dataflow_pipe_b = _RAND_1921[0:0];
  _RAND_1922 = {1{`RANDOM}};
  mesh_0_4_io_in_control_0_propagate_pipe_b = _RAND_1922[0:0];
  _RAND_1923 = {1{`RANDOM}};
  mesh_0_4_io_in_control_1_shift_pipe_b = _RAND_1923[4:0];
  _RAND_1924 = {1{`RANDOM}};
  mesh_0_4_io_in_control_1_dataflow_pipe_b = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  mesh_0_4_io_in_control_1_propagate_pipe_b = _RAND_1925[0:0];
  _RAND_1926 = {1{`RANDOM}};
  mesh_1_4_io_in_control_0_shift_pipe_b = _RAND_1926[4:0];
  _RAND_1927 = {1{`RANDOM}};
  mesh_1_4_io_in_control_0_dataflow_pipe_b = _RAND_1927[0:0];
  _RAND_1928 = {1{`RANDOM}};
  mesh_1_4_io_in_control_0_propagate_pipe_b = _RAND_1928[0:0];
  _RAND_1929 = {1{`RANDOM}};
  mesh_1_4_io_in_control_1_shift_pipe_b = _RAND_1929[4:0];
  _RAND_1930 = {1{`RANDOM}};
  mesh_1_4_io_in_control_1_dataflow_pipe_b = _RAND_1930[0:0];
  _RAND_1931 = {1{`RANDOM}};
  mesh_1_4_io_in_control_1_propagate_pipe_b = _RAND_1931[0:0];
  _RAND_1932 = {1{`RANDOM}};
  mesh_2_4_io_in_control_0_shift_pipe_b = _RAND_1932[4:0];
  _RAND_1933 = {1{`RANDOM}};
  mesh_2_4_io_in_control_0_dataflow_pipe_b = _RAND_1933[0:0];
  _RAND_1934 = {1{`RANDOM}};
  mesh_2_4_io_in_control_0_propagate_pipe_b = _RAND_1934[0:0];
  _RAND_1935 = {1{`RANDOM}};
  mesh_2_4_io_in_control_1_shift_pipe_b = _RAND_1935[4:0];
  _RAND_1936 = {1{`RANDOM}};
  mesh_2_4_io_in_control_1_dataflow_pipe_b = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  mesh_2_4_io_in_control_1_propagate_pipe_b = _RAND_1937[0:0];
  _RAND_1938 = {1{`RANDOM}};
  mesh_3_4_io_in_control_0_shift_pipe_b = _RAND_1938[4:0];
  _RAND_1939 = {1{`RANDOM}};
  mesh_3_4_io_in_control_0_dataflow_pipe_b = _RAND_1939[0:0];
  _RAND_1940 = {1{`RANDOM}};
  mesh_3_4_io_in_control_0_propagate_pipe_b = _RAND_1940[0:0];
  _RAND_1941 = {1{`RANDOM}};
  mesh_3_4_io_in_control_1_shift_pipe_b = _RAND_1941[4:0];
  _RAND_1942 = {1{`RANDOM}};
  mesh_3_4_io_in_control_1_dataflow_pipe_b = _RAND_1942[0:0];
  _RAND_1943 = {1{`RANDOM}};
  mesh_3_4_io_in_control_1_propagate_pipe_b = _RAND_1943[0:0];
  _RAND_1944 = {1{`RANDOM}};
  mesh_4_4_io_in_control_0_shift_pipe_b = _RAND_1944[4:0];
  _RAND_1945 = {1{`RANDOM}};
  mesh_4_4_io_in_control_0_dataflow_pipe_b = _RAND_1945[0:0];
  _RAND_1946 = {1{`RANDOM}};
  mesh_4_4_io_in_control_0_propagate_pipe_b = _RAND_1946[0:0];
  _RAND_1947 = {1{`RANDOM}};
  mesh_4_4_io_in_control_1_shift_pipe_b = _RAND_1947[4:0];
  _RAND_1948 = {1{`RANDOM}};
  mesh_4_4_io_in_control_1_dataflow_pipe_b = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  mesh_4_4_io_in_control_1_propagate_pipe_b = _RAND_1949[0:0];
  _RAND_1950 = {1{`RANDOM}};
  mesh_5_4_io_in_control_0_shift_pipe_b = _RAND_1950[4:0];
  _RAND_1951 = {1{`RANDOM}};
  mesh_5_4_io_in_control_0_dataflow_pipe_b = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  mesh_5_4_io_in_control_0_propagate_pipe_b = _RAND_1952[0:0];
  _RAND_1953 = {1{`RANDOM}};
  mesh_5_4_io_in_control_1_shift_pipe_b = _RAND_1953[4:0];
  _RAND_1954 = {1{`RANDOM}};
  mesh_5_4_io_in_control_1_dataflow_pipe_b = _RAND_1954[0:0];
  _RAND_1955 = {1{`RANDOM}};
  mesh_5_4_io_in_control_1_propagate_pipe_b = _RAND_1955[0:0];
  _RAND_1956 = {1{`RANDOM}};
  mesh_6_4_io_in_control_0_shift_pipe_b = _RAND_1956[4:0];
  _RAND_1957 = {1{`RANDOM}};
  mesh_6_4_io_in_control_0_dataflow_pipe_b = _RAND_1957[0:0];
  _RAND_1958 = {1{`RANDOM}};
  mesh_6_4_io_in_control_0_propagate_pipe_b = _RAND_1958[0:0];
  _RAND_1959 = {1{`RANDOM}};
  mesh_6_4_io_in_control_1_shift_pipe_b = _RAND_1959[4:0];
  _RAND_1960 = {1{`RANDOM}};
  mesh_6_4_io_in_control_1_dataflow_pipe_b = _RAND_1960[0:0];
  _RAND_1961 = {1{`RANDOM}};
  mesh_6_4_io_in_control_1_propagate_pipe_b = _RAND_1961[0:0];
  _RAND_1962 = {1{`RANDOM}};
  mesh_7_4_io_in_control_0_shift_pipe_b = _RAND_1962[4:0];
  _RAND_1963 = {1{`RANDOM}};
  mesh_7_4_io_in_control_0_dataflow_pipe_b = _RAND_1963[0:0];
  _RAND_1964 = {1{`RANDOM}};
  mesh_7_4_io_in_control_0_propagate_pipe_b = _RAND_1964[0:0];
  _RAND_1965 = {1{`RANDOM}};
  mesh_7_4_io_in_control_1_shift_pipe_b = _RAND_1965[4:0];
  _RAND_1966 = {1{`RANDOM}};
  mesh_7_4_io_in_control_1_dataflow_pipe_b = _RAND_1966[0:0];
  _RAND_1967 = {1{`RANDOM}};
  mesh_7_4_io_in_control_1_propagate_pipe_b = _RAND_1967[0:0];
  _RAND_1968 = {1{`RANDOM}};
  mesh_8_4_io_in_control_0_shift_pipe_b = _RAND_1968[4:0];
  _RAND_1969 = {1{`RANDOM}};
  mesh_8_4_io_in_control_0_dataflow_pipe_b = _RAND_1969[0:0];
  _RAND_1970 = {1{`RANDOM}};
  mesh_8_4_io_in_control_0_propagate_pipe_b = _RAND_1970[0:0];
  _RAND_1971 = {1{`RANDOM}};
  mesh_8_4_io_in_control_1_shift_pipe_b = _RAND_1971[4:0];
  _RAND_1972 = {1{`RANDOM}};
  mesh_8_4_io_in_control_1_dataflow_pipe_b = _RAND_1972[0:0];
  _RAND_1973 = {1{`RANDOM}};
  mesh_8_4_io_in_control_1_propagate_pipe_b = _RAND_1973[0:0];
  _RAND_1974 = {1{`RANDOM}};
  mesh_9_4_io_in_control_0_shift_pipe_b = _RAND_1974[4:0];
  _RAND_1975 = {1{`RANDOM}};
  mesh_9_4_io_in_control_0_dataflow_pipe_b = _RAND_1975[0:0];
  _RAND_1976 = {1{`RANDOM}};
  mesh_9_4_io_in_control_0_propagate_pipe_b = _RAND_1976[0:0];
  _RAND_1977 = {1{`RANDOM}};
  mesh_9_4_io_in_control_1_shift_pipe_b = _RAND_1977[4:0];
  _RAND_1978 = {1{`RANDOM}};
  mesh_9_4_io_in_control_1_dataflow_pipe_b = _RAND_1978[0:0];
  _RAND_1979 = {1{`RANDOM}};
  mesh_9_4_io_in_control_1_propagate_pipe_b = _RAND_1979[0:0];
  _RAND_1980 = {1{`RANDOM}};
  mesh_10_4_io_in_control_0_shift_pipe_b = _RAND_1980[4:0];
  _RAND_1981 = {1{`RANDOM}};
  mesh_10_4_io_in_control_0_dataflow_pipe_b = _RAND_1981[0:0];
  _RAND_1982 = {1{`RANDOM}};
  mesh_10_4_io_in_control_0_propagate_pipe_b = _RAND_1982[0:0];
  _RAND_1983 = {1{`RANDOM}};
  mesh_10_4_io_in_control_1_shift_pipe_b = _RAND_1983[4:0];
  _RAND_1984 = {1{`RANDOM}};
  mesh_10_4_io_in_control_1_dataflow_pipe_b = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  mesh_10_4_io_in_control_1_propagate_pipe_b = _RAND_1985[0:0];
  _RAND_1986 = {1{`RANDOM}};
  mesh_11_4_io_in_control_0_shift_pipe_b = _RAND_1986[4:0];
  _RAND_1987 = {1{`RANDOM}};
  mesh_11_4_io_in_control_0_dataflow_pipe_b = _RAND_1987[0:0];
  _RAND_1988 = {1{`RANDOM}};
  mesh_11_4_io_in_control_0_propagate_pipe_b = _RAND_1988[0:0];
  _RAND_1989 = {1{`RANDOM}};
  mesh_11_4_io_in_control_1_shift_pipe_b = _RAND_1989[4:0];
  _RAND_1990 = {1{`RANDOM}};
  mesh_11_4_io_in_control_1_dataflow_pipe_b = _RAND_1990[0:0];
  _RAND_1991 = {1{`RANDOM}};
  mesh_11_4_io_in_control_1_propagate_pipe_b = _RAND_1991[0:0];
  _RAND_1992 = {1{`RANDOM}};
  mesh_12_4_io_in_control_0_shift_pipe_b = _RAND_1992[4:0];
  _RAND_1993 = {1{`RANDOM}};
  mesh_12_4_io_in_control_0_dataflow_pipe_b = _RAND_1993[0:0];
  _RAND_1994 = {1{`RANDOM}};
  mesh_12_4_io_in_control_0_propagate_pipe_b = _RAND_1994[0:0];
  _RAND_1995 = {1{`RANDOM}};
  mesh_12_4_io_in_control_1_shift_pipe_b = _RAND_1995[4:0];
  _RAND_1996 = {1{`RANDOM}};
  mesh_12_4_io_in_control_1_dataflow_pipe_b = _RAND_1996[0:0];
  _RAND_1997 = {1{`RANDOM}};
  mesh_12_4_io_in_control_1_propagate_pipe_b = _RAND_1997[0:0];
  _RAND_1998 = {1{`RANDOM}};
  mesh_13_4_io_in_control_0_shift_pipe_b = _RAND_1998[4:0];
  _RAND_1999 = {1{`RANDOM}};
  mesh_13_4_io_in_control_0_dataflow_pipe_b = _RAND_1999[0:0];
  _RAND_2000 = {1{`RANDOM}};
  mesh_13_4_io_in_control_0_propagate_pipe_b = _RAND_2000[0:0];
  _RAND_2001 = {1{`RANDOM}};
  mesh_13_4_io_in_control_1_shift_pipe_b = _RAND_2001[4:0];
  _RAND_2002 = {1{`RANDOM}};
  mesh_13_4_io_in_control_1_dataflow_pipe_b = _RAND_2002[0:0];
  _RAND_2003 = {1{`RANDOM}};
  mesh_13_4_io_in_control_1_propagate_pipe_b = _RAND_2003[0:0];
  _RAND_2004 = {1{`RANDOM}};
  mesh_14_4_io_in_control_0_shift_pipe_b = _RAND_2004[4:0];
  _RAND_2005 = {1{`RANDOM}};
  mesh_14_4_io_in_control_0_dataflow_pipe_b = _RAND_2005[0:0];
  _RAND_2006 = {1{`RANDOM}};
  mesh_14_4_io_in_control_0_propagate_pipe_b = _RAND_2006[0:0];
  _RAND_2007 = {1{`RANDOM}};
  mesh_14_4_io_in_control_1_shift_pipe_b = _RAND_2007[4:0];
  _RAND_2008 = {1{`RANDOM}};
  mesh_14_4_io_in_control_1_dataflow_pipe_b = _RAND_2008[0:0];
  _RAND_2009 = {1{`RANDOM}};
  mesh_14_4_io_in_control_1_propagate_pipe_b = _RAND_2009[0:0];
  _RAND_2010 = {1{`RANDOM}};
  mesh_15_4_io_in_control_0_shift_pipe_b = _RAND_2010[4:0];
  _RAND_2011 = {1{`RANDOM}};
  mesh_15_4_io_in_control_0_dataflow_pipe_b = _RAND_2011[0:0];
  _RAND_2012 = {1{`RANDOM}};
  mesh_15_4_io_in_control_0_propagate_pipe_b = _RAND_2012[0:0];
  _RAND_2013 = {1{`RANDOM}};
  mesh_15_4_io_in_control_1_shift_pipe_b = _RAND_2013[4:0];
  _RAND_2014 = {1{`RANDOM}};
  mesh_15_4_io_in_control_1_dataflow_pipe_b = _RAND_2014[0:0];
  _RAND_2015 = {1{`RANDOM}};
  mesh_15_4_io_in_control_1_propagate_pipe_b = _RAND_2015[0:0];
  _RAND_2016 = {1{`RANDOM}};
  mesh_0_5_io_in_control_0_shift_pipe_b = _RAND_2016[4:0];
  _RAND_2017 = {1{`RANDOM}};
  mesh_0_5_io_in_control_0_dataflow_pipe_b = _RAND_2017[0:0];
  _RAND_2018 = {1{`RANDOM}};
  mesh_0_5_io_in_control_0_propagate_pipe_b = _RAND_2018[0:0];
  _RAND_2019 = {1{`RANDOM}};
  mesh_0_5_io_in_control_1_shift_pipe_b = _RAND_2019[4:0];
  _RAND_2020 = {1{`RANDOM}};
  mesh_0_5_io_in_control_1_dataflow_pipe_b = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  mesh_0_5_io_in_control_1_propagate_pipe_b = _RAND_2021[0:0];
  _RAND_2022 = {1{`RANDOM}};
  mesh_1_5_io_in_control_0_shift_pipe_b = _RAND_2022[4:0];
  _RAND_2023 = {1{`RANDOM}};
  mesh_1_5_io_in_control_0_dataflow_pipe_b = _RAND_2023[0:0];
  _RAND_2024 = {1{`RANDOM}};
  mesh_1_5_io_in_control_0_propagate_pipe_b = _RAND_2024[0:0];
  _RAND_2025 = {1{`RANDOM}};
  mesh_1_5_io_in_control_1_shift_pipe_b = _RAND_2025[4:0];
  _RAND_2026 = {1{`RANDOM}};
  mesh_1_5_io_in_control_1_dataflow_pipe_b = _RAND_2026[0:0];
  _RAND_2027 = {1{`RANDOM}};
  mesh_1_5_io_in_control_1_propagate_pipe_b = _RAND_2027[0:0];
  _RAND_2028 = {1{`RANDOM}};
  mesh_2_5_io_in_control_0_shift_pipe_b = _RAND_2028[4:0];
  _RAND_2029 = {1{`RANDOM}};
  mesh_2_5_io_in_control_0_dataflow_pipe_b = _RAND_2029[0:0];
  _RAND_2030 = {1{`RANDOM}};
  mesh_2_5_io_in_control_0_propagate_pipe_b = _RAND_2030[0:0];
  _RAND_2031 = {1{`RANDOM}};
  mesh_2_5_io_in_control_1_shift_pipe_b = _RAND_2031[4:0];
  _RAND_2032 = {1{`RANDOM}};
  mesh_2_5_io_in_control_1_dataflow_pipe_b = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  mesh_2_5_io_in_control_1_propagate_pipe_b = _RAND_2033[0:0];
  _RAND_2034 = {1{`RANDOM}};
  mesh_3_5_io_in_control_0_shift_pipe_b = _RAND_2034[4:0];
  _RAND_2035 = {1{`RANDOM}};
  mesh_3_5_io_in_control_0_dataflow_pipe_b = _RAND_2035[0:0];
  _RAND_2036 = {1{`RANDOM}};
  mesh_3_5_io_in_control_0_propagate_pipe_b = _RAND_2036[0:0];
  _RAND_2037 = {1{`RANDOM}};
  mesh_3_5_io_in_control_1_shift_pipe_b = _RAND_2037[4:0];
  _RAND_2038 = {1{`RANDOM}};
  mesh_3_5_io_in_control_1_dataflow_pipe_b = _RAND_2038[0:0];
  _RAND_2039 = {1{`RANDOM}};
  mesh_3_5_io_in_control_1_propagate_pipe_b = _RAND_2039[0:0];
  _RAND_2040 = {1{`RANDOM}};
  mesh_4_5_io_in_control_0_shift_pipe_b = _RAND_2040[4:0];
  _RAND_2041 = {1{`RANDOM}};
  mesh_4_5_io_in_control_0_dataflow_pipe_b = _RAND_2041[0:0];
  _RAND_2042 = {1{`RANDOM}};
  mesh_4_5_io_in_control_0_propagate_pipe_b = _RAND_2042[0:0];
  _RAND_2043 = {1{`RANDOM}};
  mesh_4_5_io_in_control_1_shift_pipe_b = _RAND_2043[4:0];
  _RAND_2044 = {1{`RANDOM}};
  mesh_4_5_io_in_control_1_dataflow_pipe_b = _RAND_2044[0:0];
  _RAND_2045 = {1{`RANDOM}};
  mesh_4_5_io_in_control_1_propagate_pipe_b = _RAND_2045[0:0];
  _RAND_2046 = {1{`RANDOM}};
  mesh_5_5_io_in_control_0_shift_pipe_b = _RAND_2046[4:0];
  _RAND_2047 = {1{`RANDOM}};
  mesh_5_5_io_in_control_0_dataflow_pipe_b = _RAND_2047[0:0];
  _RAND_2048 = {1{`RANDOM}};
  mesh_5_5_io_in_control_0_propagate_pipe_b = _RAND_2048[0:0];
  _RAND_2049 = {1{`RANDOM}};
  mesh_5_5_io_in_control_1_shift_pipe_b = _RAND_2049[4:0];
  _RAND_2050 = {1{`RANDOM}};
  mesh_5_5_io_in_control_1_dataflow_pipe_b = _RAND_2050[0:0];
  _RAND_2051 = {1{`RANDOM}};
  mesh_5_5_io_in_control_1_propagate_pipe_b = _RAND_2051[0:0];
  _RAND_2052 = {1{`RANDOM}};
  mesh_6_5_io_in_control_0_shift_pipe_b = _RAND_2052[4:0];
  _RAND_2053 = {1{`RANDOM}};
  mesh_6_5_io_in_control_0_dataflow_pipe_b = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  mesh_6_5_io_in_control_0_propagate_pipe_b = _RAND_2054[0:0];
  _RAND_2055 = {1{`RANDOM}};
  mesh_6_5_io_in_control_1_shift_pipe_b = _RAND_2055[4:0];
  _RAND_2056 = {1{`RANDOM}};
  mesh_6_5_io_in_control_1_dataflow_pipe_b = _RAND_2056[0:0];
  _RAND_2057 = {1{`RANDOM}};
  mesh_6_5_io_in_control_1_propagate_pipe_b = _RAND_2057[0:0];
  _RAND_2058 = {1{`RANDOM}};
  mesh_7_5_io_in_control_0_shift_pipe_b = _RAND_2058[4:0];
  _RAND_2059 = {1{`RANDOM}};
  mesh_7_5_io_in_control_0_dataflow_pipe_b = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  mesh_7_5_io_in_control_0_propagate_pipe_b = _RAND_2060[0:0];
  _RAND_2061 = {1{`RANDOM}};
  mesh_7_5_io_in_control_1_shift_pipe_b = _RAND_2061[4:0];
  _RAND_2062 = {1{`RANDOM}};
  mesh_7_5_io_in_control_1_dataflow_pipe_b = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  mesh_7_5_io_in_control_1_propagate_pipe_b = _RAND_2063[0:0];
  _RAND_2064 = {1{`RANDOM}};
  mesh_8_5_io_in_control_0_shift_pipe_b = _RAND_2064[4:0];
  _RAND_2065 = {1{`RANDOM}};
  mesh_8_5_io_in_control_0_dataflow_pipe_b = _RAND_2065[0:0];
  _RAND_2066 = {1{`RANDOM}};
  mesh_8_5_io_in_control_0_propagate_pipe_b = _RAND_2066[0:0];
  _RAND_2067 = {1{`RANDOM}};
  mesh_8_5_io_in_control_1_shift_pipe_b = _RAND_2067[4:0];
  _RAND_2068 = {1{`RANDOM}};
  mesh_8_5_io_in_control_1_dataflow_pipe_b = _RAND_2068[0:0];
  _RAND_2069 = {1{`RANDOM}};
  mesh_8_5_io_in_control_1_propagate_pipe_b = _RAND_2069[0:0];
  _RAND_2070 = {1{`RANDOM}};
  mesh_9_5_io_in_control_0_shift_pipe_b = _RAND_2070[4:0];
  _RAND_2071 = {1{`RANDOM}};
  mesh_9_5_io_in_control_0_dataflow_pipe_b = _RAND_2071[0:0];
  _RAND_2072 = {1{`RANDOM}};
  mesh_9_5_io_in_control_0_propagate_pipe_b = _RAND_2072[0:0];
  _RAND_2073 = {1{`RANDOM}};
  mesh_9_5_io_in_control_1_shift_pipe_b = _RAND_2073[4:0];
  _RAND_2074 = {1{`RANDOM}};
  mesh_9_5_io_in_control_1_dataflow_pipe_b = _RAND_2074[0:0];
  _RAND_2075 = {1{`RANDOM}};
  mesh_9_5_io_in_control_1_propagate_pipe_b = _RAND_2075[0:0];
  _RAND_2076 = {1{`RANDOM}};
  mesh_10_5_io_in_control_0_shift_pipe_b = _RAND_2076[4:0];
  _RAND_2077 = {1{`RANDOM}};
  mesh_10_5_io_in_control_0_dataflow_pipe_b = _RAND_2077[0:0];
  _RAND_2078 = {1{`RANDOM}};
  mesh_10_5_io_in_control_0_propagate_pipe_b = _RAND_2078[0:0];
  _RAND_2079 = {1{`RANDOM}};
  mesh_10_5_io_in_control_1_shift_pipe_b = _RAND_2079[4:0];
  _RAND_2080 = {1{`RANDOM}};
  mesh_10_5_io_in_control_1_dataflow_pipe_b = _RAND_2080[0:0];
  _RAND_2081 = {1{`RANDOM}};
  mesh_10_5_io_in_control_1_propagate_pipe_b = _RAND_2081[0:0];
  _RAND_2082 = {1{`RANDOM}};
  mesh_11_5_io_in_control_0_shift_pipe_b = _RAND_2082[4:0];
  _RAND_2083 = {1{`RANDOM}};
  mesh_11_5_io_in_control_0_dataflow_pipe_b = _RAND_2083[0:0];
  _RAND_2084 = {1{`RANDOM}};
  mesh_11_5_io_in_control_0_propagate_pipe_b = _RAND_2084[0:0];
  _RAND_2085 = {1{`RANDOM}};
  mesh_11_5_io_in_control_1_shift_pipe_b = _RAND_2085[4:0];
  _RAND_2086 = {1{`RANDOM}};
  mesh_11_5_io_in_control_1_dataflow_pipe_b = _RAND_2086[0:0];
  _RAND_2087 = {1{`RANDOM}};
  mesh_11_5_io_in_control_1_propagate_pipe_b = _RAND_2087[0:0];
  _RAND_2088 = {1{`RANDOM}};
  mesh_12_5_io_in_control_0_shift_pipe_b = _RAND_2088[4:0];
  _RAND_2089 = {1{`RANDOM}};
  mesh_12_5_io_in_control_0_dataflow_pipe_b = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  mesh_12_5_io_in_control_0_propagate_pipe_b = _RAND_2090[0:0];
  _RAND_2091 = {1{`RANDOM}};
  mesh_12_5_io_in_control_1_shift_pipe_b = _RAND_2091[4:0];
  _RAND_2092 = {1{`RANDOM}};
  mesh_12_5_io_in_control_1_dataflow_pipe_b = _RAND_2092[0:0];
  _RAND_2093 = {1{`RANDOM}};
  mesh_12_5_io_in_control_1_propagate_pipe_b = _RAND_2093[0:0];
  _RAND_2094 = {1{`RANDOM}};
  mesh_13_5_io_in_control_0_shift_pipe_b = _RAND_2094[4:0];
  _RAND_2095 = {1{`RANDOM}};
  mesh_13_5_io_in_control_0_dataflow_pipe_b = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  mesh_13_5_io_in_control_0_propagate_pipe_b = _RAND_2096[0:0];
  _RAND_2097 = {1{`RANDOM}};
  mesh_13_5_io_in_control_1_shift_pipe_b = _RAND_2097[4:0];
  _RAND_2098 = {1{`RANDOM}};
  mesh_13_5_io_in_control_1_dataflow_pipe_b = _RAND_2098[0:0];
  _RAND_2099 = {1{`RANDOM}};
  mesh_13_5_io_in_control_1_propagate_pipe_b = _RAND_2099[0:0];
  _RAND_2100 = {1{`RANDOM}};
  mesh_14_5_io_in_control_0_shift_pipe_b = _RAND_2100[4:0];
  _RAND_2101 = {1{`RANDOM}};
  mesh_14_5_io_in_control_0_dataflow_pipe_b = _RAND_2101[0:0];
  _RAND_2102 = {1{`RANDOM}};
  mesh_14_5_io_in_control_0_propagate_pipe_b = _RAND_2102[0:0];
  _RAND_2103 = {1{`RANDOM}};
  mesh_14_5_io_in_control_1_shift_pipe_b = _RAND_2103[4:0];
  _RAND_2104 = {1{`RANDOM}};
  mesh_14_5_io_in_control_1_dataflow_pipe_b = _RAND_2104[0:0];
  _RAND_2105 = {1{`RANDOM}};
  mesh_14_5_io_in_control_1_propagate_pipe_b = _RAND_2105[0:0];
  _RAND_2106 = {1{`RANDOM}};
  mesh_15_5_io_in_control_0_shift_pipe_b = _RAND_2106[4:0];
  _RAND_2107 = {1{`RANDOM}};
  mesh_15_5_io_in_control_0_dataflow_pipe_b = _RAND_2107[0:0];
  _RAND_2108 = {1{`RANDOM}};
  mesh_15_5_io_in_control_0_propagate_pipe_b = _RAND_2108[0:0];
  _RAND_2109 = {1{`RANDOM}};
  mesh_15_5_io_in_control_1_shift_pipe_b = _RAND_2109[4:0];
  _RAND_2110 = {1{`RANDOM}};
  mesh_15_5_io_in_control_1_dataflow_pipe_b = _RAND_2110[0:0];
  _RAND_2111 = {1{`RANDOM}};
  mesh_15_5_io_in_control_1_propagate_pipe_b = _RAND_2111[0:0];
  _RAND_2112 = {1{`RANDOM}};
  mesh_0_6_io_in_control_0_shift_pipe_b = _RAND_2112[4:0];
  _RAND_2113 = {1{`RANDOM}};
  mesh_0_6_io_in_control_0_dataflow_pipe_b = _RAND_2113[0:0];
  _RAND_2114 = {1{`RANDOM}};
  mesh_0_6_io_in_control_0_propagate_pipe_b = _RAND_2114[0:0];
  _RAND_2115 = {1{`RANDOM}};
  mesh_0_6_io_in_control_1_shift_pipe_b = _RAND_2115[4:0];
  _RAND_2116 = {1{`RANDOM}};
  mesh_0_6_io_in_control_1_dataflow_pipe_b = _RAND_2116[0:0];
  _RAND_2117 = {1{`RANDOM}};
  mesh_0_6_io_in_control_1_propagate_pipe_b = _RAND_2117[0:0];
  _RAND_2118 = {1{`RANDOM}};
  mesh_1_6_io_in_control_0_shift_pipe_b = _RAND_2118[4:0];
  _RAND_2119 = {1{`RANDOM}};
  mesh_1_6_io_in_control_0_dataflow_pipe_b = _RAND_2119[0:0];
  _RAND_2120 = {1{`RANDOM}};
  mesh_1_6_io_in_control_0_propagate_pipe_b = _RAND_2120[0:0];
  _RAND_2121 = {1{`RANDOM}};
  mesh_1_6_io_in_control_1_shift_pipe_b = _RAND_2121[4:0];
  _RAND_2122 = {1{`RANDOM}};
  mesh_1_6_io_in_control_1_dataflow_pipe_b = _RAND_2122[0:0];
  _RAND_2123 = {1{`RANDOM}};
  mesh_1_6_io_in_control_1_propagate_pipe_b = _RAND_2123[0:0];
  _RAND_2124 = {1{`RANDOM}};
  mesh_2_6_io_in_control_0_shift_pipe_b = _RAND_2124[4:0];
  _RAND_2125 = {1{`RANDOM}};
  mesh_2_6_io_in_control_0_dataflow_pipe_b = _RAND_2125[0:0];
  _RAND_2126 = {1{`RANDOM}};
  mesh_2_6_io_in_control_0_propagate_pipe_b = _RAND_2126[0:0];
  _RAND_2127 = {1{`RANDOM}};
  mesh_2_6_io_in_control_1_shift_pipe_b = _RAND_2127[4:0];
  _RAND_2128 = {1{`RANDOM}};
  mesh_2_6_io_in_control_1_dataflow_pipe_b = _RAND_2128[0:0];
  _RAND_2129 = {1{`RANDOM}};
  mesh_2_6_io_in_control_1_propagate_pipe_b = _RAND_2129[0:0];
  _RAND_2130 = {1{`RANDOM}};
  mesh_3_6_io_in_control_0_shift_pipe_b = _RAND_2130[4:0];
  _RAND_2131 = {1{`RANDOM}};
  mesh_3_6_io_in_control_0_dataflow_pipe_b = _RAND_2131[0:0];
  _RAND_2132 = {1{`RANDOM}};
  mesh_3_6_io_in_control_0_propagate_pipe_b = _RAND_2132[0:0];
  _RAND_2133 = {1{`RANDOM}};
  mesh_3_6_io_in_control_1_shift_pipe_b = _RAND_2133[4:0];
  _RAND_2134 = {1{`RANDOM}};
  mesh_3_6_io_in_control_1_dataflow_pipe_b = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  mesh_3_6_io_in_control_1_propagate_pipe_b = _RAND_2135[0:0];
  _RAND_2136 = {1{`RANDOM}};
  mesh_4_6_io_in_control_0_shift_pipe_b = _RAND_2136[4:0];
  _RAND_2137 = {1{`RANDOM}};
  mesh_4_6_io_in_control_0_dataflow_pipe_b = _RAND_2137[0:0];
  _RAND_2138 = {1{`RANDOM}};
  mesh_4_6_io_in_control_0_propagate_pipe_b = _RAND_2138[0:0];
  _RAND_2139 = {1{`RANDOM}};
  mesh_4_6_io_in_control_1_shift_pipe_b = _RAND_2139[4:0];
  _RAND_2140 = {1{`RANDOM}};
  mesh_4_6_io_in_control_1_dataflow_pipe_b = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  mesh_4_6_io_in_control_1_propagate_pipe_b = _RAND_2141[0:0];
  _RAND_2142 = {1{`RANDOM}};
  mesh_5_6_io_in_control_0_shift_pipe_b = _RAND_2142[4:0];
  _RAND_2143 = {1{`RANDOM}};
  mesh_5_6_io_in_control_0_dataflow_pipe_b = _RAND_2143[0:0];
  _RAND_2144 = {1{`RANDOM}};
  mesh_5_6_io_in_control_0_propagate_pipe_b = _RAND_2144[0:0];
  _RAND_2145 = {1{`RANDOM}};
  mesh_5_6_io_in_control_1_shift_pipe_b = _RAND_2145[4:0];
  _RAND_2146 = {1{`RANDOM}};
  mesh_5_6_io_in_control_1_dataflow_pipe_b = _RAND_2146[0:0];
  _RAND_2147 = {1{`RANDOM}};
  mesh_5_6_io_in_control_1_propagate_pipe_b = _RAND_2147[0:0];
  _RAND_2148 = {1{`RANDOM}};
  mesh_6_6_io_in_control_0_shift_pipe_b = _RAND_2148[4:0];
  _RAND_2149 = {1{`RANDOM}};
  mesh_6_6_io_in_control_0_dataflow_pipe_b = _RAND_2149[0:0];
  _RAND_2150 = {1{`RANDOM}};
  mesh_6_6_io_in_control_0_propagate_pipe_b = _RAND_2150[0:0];
  _RAND_2151 = {1{`RANDOM}};
  mesh_6_6_io_in_control_1_shift_pipe_b = _RAND_2151[4:0];
  _RAND_2152 = {1{`RANDOM}};
  mesh_6_6_io_in_control_1_dataflow_pipe_b = _RAND_2152[0:0];
  _RAND_2153 = {1{`RANDOM}};
  mesh_6_6_io_in_control_1_propagate_pipe_b = _RAND_2153[0:0];
  _RAND_2154 = {1{`RANDOM}};
  mesh_7_6_io_in_control_0_shift_pipe_b = _RAND_2154[4:0];
  _RAND_2155 = {1{`RANDOM}};
  mesh_7_6_io_in_control_0_dataflow_pipe_b = _RAND_2155[0:0];
  _RAND_2156 = {1{`RANDOM}};
  mesh_7_6_io_in_control_0_propagate_pipe_b = _RAND_2156[0:0];
  _RAND_2157 = {1{`RANDOM}};
  mesh_7_6_io_in_control_1_shift_pipe_b = _RAND_2157[4:0];
  _RAND_2158 = {1{`RANDOM}};
  mesh_7_6_io_in_control_1_dataflow_pipe_b = _RAND_2158[0:0];
  _RAND_2159 = {1{`RANDOM}};
  mesh_7_6_io_in_control_1_propagate_pipe_b = _RAND_2159[0:0];
  _RAND_2160 = {1{`RANDOM}};
  mesh_8_6_io_in_control_0_shift_pipe_b = _RAND_2160[4:0];
  _RAND_2161 = {1{`RANDOM}};
  mesh_8_6_io_in_control_0_dataflow_pipe_b = _RAND_2161[0:0];
  _RAND_2162 = {1{`RANDOM}};
  mesh_8_6_io_in_control_0_propagate_pipe_b = _RAND_2162[0:0];
  _RAND_2163 = {1{`RANDOM}};
  mesh_8_6_io_in_control_1_shift_pipe_b = _RAND_2163[4:0];
  _RAND_2164 = {1{`RANDOM}};
  mesh_8_6_io_in_control_1_dataflow_pipe_b = _RAND_2164[0:0];
  _RAND_2165 = {1{`RANDOM}};
  mesh_8_6_io_in_control_1_propagate_pipe_b = _RAND_2165[0:0];
  _RAND_2166 = {1{`RANDOM}};
  mesh_9_6_io_in_control_0_shift_pipe_b = _RAND_2166[4:0];
  _RAND_2167 = {1{`RANDOM}};
  mesh_9_6_io_in_control_0_dataflow_pipe_b = _RAND_2167[0:0];
  _RAND_2168 = {1{`RANDOM}};
  mesh_9_6_io_in_control_0_propagate_pipe_b = _RAND_2168[0:0];
  _RAND_2169 = {1{`RANDOM}};
  mesh_9_6_io_in_control_1_shift_pipe_b = _RAND_2169[4:0];
  _RAND_2170 = {1{`RANDOM}};
  mesh_9_6_io_in_control_1_dataflow_pipe_b = _RAND_2170[0:0];
  _RAND_2171 = {1{`RANDOM}};
  mesh_9_6_io_in_control_1_propagate_pipe_b = _RAND_2171[0:0];
  _RAND_2172 = {1{`RANDOM}};
  mesh_10_6_io_in_control_0_shift_pipe_b = _RAND_2172[4:0];
  _RAND_2173 = {1{`RANDOM}};
  mesh_10_6_io_in_control_0_dataflow_pipe_b = _RAND_2173[0:0];
  _RAND_2174 = {1{`RANDOM}};
  mesh_10_6_io_in_control_0_propagate_pipe_b = _RAND_2174[0:0];
  _RAND_2175 = {1{`RANDOM}};
  mesh_10_6_io_in_control_1_shift_pipe_b = _RAND_2175[4:0];
  _RAND_2176 = {1{`RANDOM}};
  mesh_10_6_io_in_control_1_dataflow_pipe_b = _RAND_2176[0:0];
  _RAND_2177 = {1{`RANDOM}};
  mesh_10_6_io_in_control_1_propagate_pipe_b = _RAND_2177[0:0];
  _RAND_2178 = {1{`RANDOM}};
  mesh_11_6_io_in_control_0_shift_pipe_b = _RAND_2178[4:0];
  _RAND_2179 = {1{`RANDOM}};
  mesh_11_6_io_in_control_0_dataflow_pipe_b = _RAND_2179[0:0];
  _RAND_2180 = {1{`RANDOM}};
  mesh_11_6_io_in_control_0_propagate_pipe_b = _RAND_2180[0:0];
  _RAND_2181 = {1{`RANDOM}};
  mesh_11_6_io_in_control_1_shift_pipe_b = _RAND_2181[4:0];
  _RAND_2182 = {1{`RANDOM}};
  mesh_11_6_io_in_control_1_dataflow_pipe_b = _RAND_2182[0:0];
  _RAND_2183 = {1{`RANDOM}};
  mesh_11_6_io_in_control_1_propagate_pipe_b = _RAND_2183[0:0];
  _RAND_2184 = {1{`RANDOM}};
  mesh_12_6_io_in_control_0_shift_pipe_b = _RAND_2184[4:0];
  _RAND_2185 = {1{`RANDOM}};
  mesh_12_6_io_in_control_0_dataflow_pipe_b = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  mesh_12_6_io_in_control_0_propagate_pipe_b = _RAND_2186[0:0];
  _RAND_2187 = {1{`RANDOM}};
  mesh_12_6_io_in_control_1_shift_pipe_b = _RAND_2187[4:0];
  _RAND_2188 = {1{`RANDOM}};
  mesh_12_6_io_in_control_1_dataflow_pipe_b = _RAND_2188[0:0];
  _RAND_2189 = {1{`RANDOM}};
  mesh_12_6_io_in_control_1_propagate_pipe_b = _RAND_2189[0:0];
  _RAND_2190 = {1{`RANDOM}};
  mesh_13_6_io_in_control_0_shift_pipe_b = _RAND_2190[4:0];
  _RAND_2191 = {1{`RANDOM}};
  mesh_13_6_io_in_control_0_dataflow_pipe_b = _RAND_2191[0:0];
  _RAND_2192 = {1{`RANDOM}};
  mesh_13_6_io_in_control_0_propagate_pipe_b = _RAND_2192[0:0];
  _RAND_2193 = {1{`RANDOM}};
  mesh_13_6_io_in_control_1_shift_pipe_b = _RAND_2193[4:0];
  _RAND_2194 = {1{`RANDOM}};
  mesh_13_6_io_in_control_1_dataflow_pipe_b = _RAND_2194[0:0];
  _RAND_2195 = {1{`RANDOM}};
  mesh_13_6_io_in_control_1_propagate_pipe_b = _RAND_2195[0:0];
  _RAND_2196 = {1{`RANDOM}};
  mesh_14_6_io_in_control_0_shift_pipe_b = _RAND_2196[4:0];
  _RAND_2197 = {1{`RANDOM}};
  mesh_14_6_io_in_control_0_dataflow_pipe_b = _RAND_2197[0:0];
  _RAND_2198 = {1{`RANDOM}};
  mesh_14_6_io_in_control_0_propagate_pipe_b = _RAND_2198[0:0];
  _RAND_2199 = {1{`RANDOM}};
  mesh_14_6_io_in_control_1_shift_pipe_b = _RAND_2199[4:0];
  _RAND_2200 = {1{`RANDOM}};
  mesh_14_6_io_in_control_1_dataflow_pipe_b = _RAND_2200[0:0];
  _RAND_2201 = {1{`RANDOM}};
  mesh_14_6_io_in_control_1_propagate_pipe_b = _RAND_2201[0:0];
  _RAND_2202 = {1{`RANDOM}};
  mesh_15_6_io_in_control_0_shift_pipe_b = _RAND_2202[4:0];
  _RAND_2203 = {1{`RANDOM}};
  mesh_15_6_io_in_control_0_dataflow_pipe_b = _RAND_2203[0:0];
  _RAND_2204 = {1{`RANDOM}};
  mesh_15_6_io_in_control_0_propagate_pipe_b = _RAND_2204[0:0];
  _RAND_2205 = {1{`RANDOM}};
  mesh_15_6_io_in_control_1_shift_pipe_b = _RAND_2205[4:0];
  _RAND_2206 = {1{`RANDOM}};
  mesh_15_6_io_in_control_1_dataflow_pipe_b = _RAND_2206[0:0];
  _RAND_2207 = {1{`RANDOM}};
  mesh_15_6_io_in_control_1_propagate_pipe_b = _RAND_2207[0:0];
  _RAND_2208 = {1{`RANDOM}};
  mesh_0_7_io_in_control_0_shift_pipe_b = _RAND_2208[4:0];
  _RAND_2209 = {1{`RANDOM}};
  mesh_0_7_io_in_control_0_dataflow_pipe_b = _RAND_2209[0:0];
  _RAND_2210 = {1{`RANDOM}};
  mesh_0_7_io_in_control_0_propagate_pipe_b = _RAND_2210[0:0];
  _RAND_2211 = {1{`RANDOM}};
  mesh_0_7_io_in_control_1_shift_pipe_b = _RAND_2211[4:0];
  _RAND_2212 = {1{`RANDOM}};
  mesh_0_7_io_in_control_1_dataflow_pipe_b = _RAND_2212[0:0];
  _RAND_2213 = {1{`RANDOM}};
  mesh_0_7_io_in_control_1_propagate_pipe_b = _RAND_2213[0:0];
  _RAND_2214 = {1{`RANDOM}};
  mesh_1_7_io_in_control_0_shift_pipe_b = _RAND_2214[4:0];
  _RAND_2215 = {1{`RANDOM}};
  mesh_1_7_io_in_control_0_dataflow_pipe_b = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  mesh_1_7_io_in_control_0_propagate_pipe_b = _RAND_2216[0:0];
  _RAND_2217 = {1{`RANDOM}};
  mesh_1_7_io_in_control_1_shift_pipe_b = _RAND_2217[4:0];
  _RAND_2218 = {1{`RANDOM}};
  mesh_1_7_io_in_control_1_dataflow_pipe_b = _RAND_2218[0:0];
  _RAND_2219 = {1{`RANDOM}};
  mesh_1_7_io_in_control_1_propagate_pipe_b = _RAND_2219[0:0];
  _RAND_2220 = {1{`RANDOM}};
  mesh_2_7_io_in_control_0_shift_pipe_b = _RAND_2220[4:0];
  _RAND_2221 = {1{`RANDOM}};
  mesh_2_7_io_in_control_0_dataflow_pipe_b = _RAND_2221[0:0];
  _RAND_2222 = {1{`RANDOM}};
  mesh_2_7_io_in_control_0_propagate_pipe_b = _RAND_2222[0:0];
  _RAND_2223 = {1{`RANDOM}};
  mesh_2_7_io_in_control_1_shift_pipe_b = _RAND_2223[4:0];
  _RAND_2224 = {1{`RANDOM}};
  mesh_2_7_io_in_control_1_dataflow_pipe_b = _RAND_2224[0:0];
  _RAND_2225 = {1{`RANDOM}};
  mesh_2_7_io_in_control_1_propagate_pipe_b = _RAND_2225[0:0];
  _RAND_2226 = {1{`RANDOM}};
  mesh_3_7_io_in_control_0_shift_pipe_b = _RAND_2226[4:0];
  _RAND_2227 = {1{`RANDOM}};
  mesh_3_7_io_in_control_0_dataflow_pipe_b = _RAND_2227[0:0];
  _RAND_2228 = {1{`RANDOM}};
  mesh_3_7_io_in_control_0_propagate_pipe_b = _RAND_2228[0:0];
  _RAND_2229 = {1{`RANDOM}};
  mesh_3_7_io_in_control_1_shift_pipe_b = _RAND_2229[4:0];
  _RAND_2230 = {1{`RANDOM}};
  mesh_3_7_io_in_control_1_dataflow_pipe_b = _RAND_2230[0:0];
  _RAND_2231 = {1{`RANDOM}};
  mesh_3_7_io_in_control_1_propagate_pipe_b = _RAND_2231[0:0];
  _RAND_2232 = {1{`RANDOM}};
  mesh_4_7_io_in_control_0_shift_pipe_b = _RAND_2232[4:0];
  _RAND_2233 = {1{`RANDOM}};
  mesh_4_7_io_in_control_0_dataflow_pipe_b = _RAND_2233[0:0];
  _RAND_2234 = {1{`RANDOM}};
  mesh_4_7_io_in_control_0_propagate_pipe_b = _RAND_2234[0:0];
  _RAND_2235 = {1{`RANDOM}};
  mesh_4_7_io_in_control_1_shift_pipe_b = _RAND_2235[4:0];
  _RAND_2236 = {1{`RANDOM}};
  mesh_4_7_io_in_control_1_dataflow_pipe_b = _RAND_2236[0:0];
  _RAND_2237 = {1{`RANDOM}};
  mesh_4_7_io_in_control_1_propagate_pipe_b = _RAND_2237[0:0];
  _RAND_2238 = {1{`RANDOM}};
  mesh_5_7_io_in_control_0_shift_pipe_b = _RAND_2238[4:0];
  _RAND_2239 = {1{`RANDOM}};
  mesh_5_7_io_in_control_0_dataflow_pipe_b = _RAND_2239[0:0];
  _RAND_2240 = {1{`RANDOM}};
  mesh_5_7_io_in_control_0_propagate_pipe_b = _RAND_2240[0:0];
  _RAND_2241 = {1{`RANDOM}};
  mesh_5_7_io_in_control_1_shift_pipe_b = _RAND_2241[4:0];
  _RAND_2242 = {1{`RANDOM}};
  mesh_5_7_io_in_control_1_dataflow_pipe_b = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  mesh_5_7_io_in_control_1_propagate_pipe_b = _RAND_2243[0:0];
  _RAND_2244 = {1{`RANDOM}};
  mesh_6_7_io_in_control_0_shift_pipe_b = _RAND_2244[4:0];
  _RAND_2245 = {1{`RANDOM}};
  mesh_6_7_io_in_control_0_dataflow_pipe_b = _RAND_2245[0:0];
  _RAND_2246 = {1{`RANDOM}};
  mesh_6_7_io_in_control_0_propagate_pipe_b = _RAND_2246[0:0];
  _RAND_2247 = {1{`RANDOM}};
  mesh_6_7_io_in_control_1_shift_pipe_b = _RAND_2247[4:0];
  _RAND_2248 = {1{`RANDOM}};
  mesh_6_7_io_in_control_1_dataflow_pipe_b = _RAND_2248[0:0];
  _RAND_2249 = {1{`RANDOM}};
  mesh_6_7_io_in_control_1_propagate_pipe_b = _RAND_2249[0:0];
  _RAND_2250 = {1{`RANDOM}};
  mesh_7_7_io_in_control_0_shift_pipe_b = _RAND_2250[4:0];
  _RAND_2251 = {1{`RANDOM}};
  mesh_7_7_io_in_control_0_dataflow_pipe_b = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  mesh_7_7_io_in_control_0_propagate_pipe_b = _RAND_2252[0:0];
  _RAND_2253 = {1{`RANDOM}};
  mesh_7_7_io_in_control_1_shift_pipe_b = _RAND_2253[4:0];
  _RAND_2254 = {1{`RANDOM}};
  mesh_7_7_io_in_control_1_dataflow_pipe_b = _RAND_2254[0:0];
  _RAND_2255 = {1{`RANDOM}};
  mesh_7_7_io_in_control_1_propagate_pipe_b = _RAND_2255[0:0];
  _RAND_2256 = {1{`RANDOM}};
  mesh_8_7_io_in_control_0_shift_pipe_b = _RAND_2256[4:0];
  _RAND_2257 = {1{`RANDOM}};
  mesh_8_7_io_in_control_0_dataflow_pipe_b = _RAND_2257[0:0];
  _RAND_2258 = {1{`RANDOM}};
  mesh_8_7_io_in_control_0_propagate_pipe_b = _RAND_2258[0:0];
  _RAND_2259 = {1{`RANDOM}};
  mesh_8_7_io_in_control_1_shift_pipe_b = _RAND_2259[4:0];
  _RAND_2260 = {1{`RANDOM}};
  mesh_8_7_io_in_control_1_dataflow_pipe_b = _RAND_2260[0:0];
  _RAND_2261 = {1{`RANDOM}};
  mesh_8_7_io_in_control_1_propagate_pipe_b = _RAND_2261[0:0];
  _RAND_2262 = {1{`RANDOM}};
  mesh_9_7_io_in_control_0_shift_pipe_b = _RAND_2262[4:0];
  _RAND_2263 = {1{`RANDOM}};
  mesh_9_7_io_in_control_0_dataflow_pipe_b = _RAND_2263[0:0];
  _RAND_2264 = {1{`RANDOM}};
  mesh_9_7_io_in_control_0_propagate_pipe_b = _RAND_2264[0:0];
  _RAND_2265 = {1{`RANDOM}};
  mesh_9_7_io_in_control_1_shift_pipe_b = _RAND_2265[4:0];
  _RAND_2266 = {1{`RANDOM}};
  mesh_9_7_io_in_control_1_dataflow_pipe_b = _RAND_2266[0:0];
  _RAND_2267 = {1{`RANDOM}};
  mesh_9_7_io_in_control_1_propagate_pipe_b = _RAND_2267[0:0];
  _RAND_2268 = {1{`RANDOM}};
  mesh_10_7_io_in_control_0_shift_pipe_b = _RAND_2268[4:0];
  _RAND_2269 = {1{`RANDOM}};
  mesh_10_7_io_in_control_0_dataflow_pipe_b = _RAND_2269[0:0];
  _RAND_2270 = {1{`RANDOM}};
  mesh_10_7_io_in_control_0_propagate_pipe_b = _RAND_2270[0:0];
  _RAND_2271 = {1{`RANDOM}};
  mesh_10_7_io_in_control_1_shift_pipe_b = _RAND_2271[4:0];
  _RAND_2272 = {1{`RANDOM}};
  mesh_10_7_io_in_control_1_dataflow_pipe_b = _RAND_2272[0:0];
  _RAND_2273 = {1{`RANDOM}};
  mesh_10_7_io_in_control_1_propagate_pipe_b = _RAND_2273[0:0];
  _RAND_2274 = {1{`RANDOM}};
  mesh_11_7_io_in_control_0_shift_pipe_b = _RAND_2274[4:0];
  _RAND_2275 = {1{`RANDOM}};
  mesh_11_7_io_in_control_0_dataflow_pipe_b = _RAND_2275[0:0];
  _RAND_2276 = {1{`RANDOM}};
  mesh_11_7_io_in_control_0_propagate_pipe_b = _RAND_2276[0:0];
  _RAND_2277 = {1{`RANDOM}};
  mesh_11_7_io_in_control_1_shift_pipe_b = _RAND_2277[4:0];
  _RAND_2278 = {1{`RANDOM}};
  mesh_11_7_io_in_control_1_dataflow_pipe_b = _RAND_2278[0:0];
  _RAND_2279 = {1{`RANDOM}};
  mesh_11_7_io_in_control_1_propagate_pipe_b = _RAND_2279[0:0];
  _RAND_2280 = {1{`RANDOM}};
  mesh_12_7_io_in_control_0_shift_pipe_b = _RAND_2280[4:0];
  _RAND_2281 = {1{`RANDOM}};
  mesh_12_7_io_in_control_0_dataflow_pipe_b = _RAND_2281[0:0];
  _RAND_2282 = {1{`RANDOM}};
  mesh_12_7_io_in_control_0_propagate_pipe_b = _RAND_2282[0:0];
  _RAND_2283 = {1{`RANDOM}};
  mesh_12_7_io_in_control_1_shift_pipe_b = _RAND_2283[4:0];
  _RAND_2284 = {1{`RANDOM}};
  mesh_12_7_io_in_control_1_dataflow_pipe_b = _RAND_2284[0:0];
  _RAND_2285 = {1{`RANDOM}};
  mesh_12_7_io_in_control_1_propagate_pipe_b = _RAND_2285[0:0];
  _RAND_2286 = {1{`RANDOM}};
  mesh_13_7_io_in_control_0_shift_pipe_b = _RAND_2286[4:0];
  _RAND_2287 = {1{`RANDOM}};
  mesh_13_7_io_in_control_0_dataflow_pipe_b = _RAND_2287[0:0];
  _RAND_2288 = {1{`RANDOM}};
  mesh_13_7_io_in_control_0_propagate_pipe_b = _RAND_2288[0:0];
  _RAND_2289 = {1{`RANDOM}};
  mesh_13_7_io_in_control_1_shift_pipe_b = _RAND_2289[4:0];
  _RAND_2290 = {1{`RANDOM}};
  mesh_13_7_io_in_control_1_dataflow_pipe_b = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  mesh_13_7_io_in_control_1_propagate_pipe_b = _RAND_2291[0:0];
  _RAND_2292 = {1{`RANDOM}};
  mesh_14_7_io_in_control_0_shift_pipe_b = _RAND_2292[4:0];
  _RAND_2293 = {1{`RANDOM}};
  mesh_14_7_io_in_control_0_dataflow_pipe_b = _RAND_2293[0:0];
  _RAND_2294 = {1{`RANDOM}};
  mesh_14_7_io_in_control_0_propagate_pipe_b = _RAND_2294[0:0];
  _RAND_2295 = {1{`RANDOM}};
  mesh_14_7_io_in_control_1_shift_pipe_b = _RAND_2295[4:0];
  _RAND_2296 = {1{`RANDOM}};
  mesh_14_7_io_in_control_1_dataflow_pipe_b = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  mesh_14_7_io_in_control_1_propagate_pipe_b = _RAND_2297[0:0];
  _RAND_2298 = {1{`RANDOM}};
  mesh_15_7_io_in_control_0_shift_pipe_b = _RAND_2298[4:0];
  _RAND_2299 = {1{`RANDOM}};
  mesh_15_7_io_in_control_0_dataflow_pipe_b = _RAND_2299[0:0];
  _RAND_2300 = {1{`RANDOM}};
  mesh_15_7_io_in_control_0_propagate_pipe_b = _RAND_2300[0:0];
  _RAND_2301 = {1{`RANDOM}};
  mesh_15_7_io_in_control_1_shift_pipe_b = _RAND_2301[4:0];
  _RAND_2302 = {1{`RANDOM}};
  mesh_15_7_io_in_control_1_dataflow_pipe_b = _RAND_2302[0:0];
  _RAND_2303 = {1{`RANDOM}};
  mesh_15_7_io_in_control_1_propagate_pipe_b = _RAND_2303[0:0];
  _RAND_2304 = {1{`RANDOM}};
  mesh_0_8_io_in_control_0_shift_pipe_b = _RAND_2304[4:0];
  _RAND_2305 = {1{`RANDOM}};
  mesh_0_8_io_in_control_0_dataflow_pipe_b = _RAND_2305[0:0];
  _RAND_2306 = {1{`RANDOM}};
  mesh_0_8_io_in_control_0_propagate_pipe_b = _RAND_2306[0:0];
  _RAND_2307 = {1{`RANDOM}};
  mesh_0_8_io_in_control_1_shift_pipe_b = _RAND_2307[4:0];
  _RAND_2308 = {1{`RANDOM}};
  mesh_0_8_io_in_control_1_dataflow_pipe_b = _RAND_2308[0:0];
  _RAND_2309 = {1{`RANDOM}};
  mesh_0_8_io_in_control_1_propagate_pipe_b = _RAND_2309[0:0];
  _RAND_2310 = {1{`RANDOM}};
  mesh_1_8_io_in_control_0_shift_pipe_b = _RAND_2310[4:0];
  _RAND_2311 = {1{`RANDOM}};
  mesh_1_8_io_in_control_0_dataflow_pipe_b = _RAND_2311[0:0];
  _RAND_2312 = {1{`RANDOM}};
  mesh_1_8_io_in_control_0_propagate_pipe_b = _RAND_2312[0:0];
  _RAND_2313 = {1{`RANDOM}};
  mesh_1_8_io_in_control_1_shift_pipe_b = _RAND_2313[4:0];
  _RAND_2314 = {1{`RANDOM}};
  mesh_1_8_io_in_control_1_dataflow_pipe_b = _RAND_2314[0:0];
  _RAND_2315 = {1{`RANDOM}};
  mesh_1_8_io_in_control_1_propagate_pipe_b = _RAND_2315[0:0];
  _RAND_2316 = {1{`RANDOM}};
  mesh_2_8_io_in_control_0_shift_pipe_b = _RAND_2316[4:0];
  _RAND_2317 = {1{`RANDOM}};
  mesh_2_8_io_in_control_0_dataflow_pipe_b = _RAND_2317[0:0];
  _RAND_2318 = {1{`RANDOM}};
  mesh_2_8_io_in_control_0_propagate_pipe_b = _RAND_2318[0:0];
  _RAND_2319 = {1{`RANDOM}};
  mesh_2_8_io_in_control_1_shift_pipe_b = _RAND_2319[4:0];
  _RAND_2320 = {1{`RANDOM}};
  mesh_2_8_io_in_control_1_dataflow_pipe_b = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  mesh_2_8_io_in_control_1_propagate_pipe_b = _RAND_2321[0:0];
  _RAND_2322 = {1{`RANDOM}};
  mesh_3_8_io_in_control_0_shift_pipe_b = _RAND_2322[4:0];
  _RAND_2323 = {1{`RANDOM}};
  mesh_3_8_io_in_control_0_dataflow_pipe_b = _RAND_2323[0:0];
  _RAND_2324 = {1{`RANDOM}};
  mesh_3_8_io_in_control_0_propagate_pipe_b = _RAND_2324[0:0];
  _RAND_2325 = {1{`RANDOM}};
  mesh_3_8_io_in_control_1_shift_pipe_b = _RAND_2325[4:0];
  _RAND_2326 = {1{`RANDOM}};
  mesh_3_8_io_in_control_1_dataflow_pipe_b = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  mesh_3_8_io_in_control_1_propagate_pipe_b = _RAND_2327[0:0];
  _RAND_2328 = {1{`RANDOM}};
  mesh_4_8_io_in_control_0_shift_pipe_b = _RAND_2328[4:0];
  _RAND_2329 = {1{`RANDOM}};
  mesh_4_8_io_in_control_0_dataflow_pipe_b = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  mesh_4_8_io_in_control_0_propagate_pipe_b = _RAND_2330[0:0];
  _RAND_2331 = {1{`RANDOM}};
  mesh_4_8_io_in_control_1_shift_pipe_b = _RAND_2331[4:0];
  _RAND_2332 = {1{`RANDOM}};
  mesh_4_8_io_in_control_1_dataflow_pipe_b = _RAND_2332[0:0];
  _RAND_2333 = {1{`RANDOM}};
  mesh_4_8_io_in_control_1_propagate_pipe_b = _RAND_2333[0:0];
  _RAND_2334 = {1{`RANDOM}};
  mesh_5_8_io_in_control_0_shift_pipe_b = _RAND_2334[4:0];
  _RAND_2335 = {1{`RANDOM}};
  mesh_5_8_io_in_control_0_dataflow_pipe_b = _RAND_2335[0:0];
  _RAND_2336 = {1{`RANDOM}};
  mesh_5_8_io_in_control_0_propagate_pipe_b = _RAND_2336[0:0];
  _RAND_2337 = {1{`RANDOM}};
  mesh_5_8_io_in_control_1_shift_pipe_b = _RAND_2337[4:0];
  _RAND_2338 = {1{`RANDOM}};
  mesh_5_8_io_in_control_1_dataflow_pipe_b = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  mesh_5_8_io_in_control_1_propagate_pipe_b = _RAND_2339[0:0];
  _RAND_2340 = {1{`RANDOM}};
  mesh_6_8_io_in_control_0_shift_pipe_b = _RAND_2340[4:0];
  _RAND_2341 = {1{`RANDOM}};
  mesh_6_8_io_in_control_0_dataflow_pipe_b = _RAND_2341[0:0];
  _RAND_2342 = {1{`RANDOM}};
  mesh_6_8_io_in_control_0_propagate_pipe_b = _RAND_2342[0:0];
  _RAND_2343 = {1{`RANDOM}};
  mesh_6_8_io_in_control_1_shift_pipe_b = _RAND_2343[4:0];
  _RAND_2344 = {1{`RANDOM}};
  mesh_6_8_io_in_control_1_dataflow_pipe_b = _RAND_2344[0:0];
  _RAND_2345 = {1{`RANDOM}};
  mesh_6_8_io_in_control_1_propagate_pipe_b = _RAND_2345[0:0];
  _RAND_2346 = {1{`RANDOM}};
  mesh_7_8_io_in_control_0_shift_pipe_b = _RAND_2346[4:0];
  _RAND_2347 = {1{`RANDOM}};
  mesh_7_8_io_in_control_0_dataflow_pipe_b = _RAND_2347[0:0];
  _RAND_2348 = {1{`RANDOM}};
  mesh_7_8_io_in_control_0_propagate_pipe_b = _RAND_2348[0:0];
  _RAND_2349 = {1{`RANDOM}};
  mesh_7_8_io_in_control_1_shift_pipe_b = _RAND_2349[4:0];
  _RAND_2350 = {1{`RANDOM}};
  mesh_7_8_io_in_control_1_dataflow_pipe_b = _RAND_2350[0:0];
  _RAND_2351 = {1{`RANDOM}};
  mesh_7_8_io_in_control_1_propagate_pipe_b = _RAND_2351[0:0];
  _RAND_2352 = {1{`RANDOM}};
  mesh_8_8_io_in_control_0_shift_pipe_b = _RAND_2352[4:0];
  _RAND_2353 = {1{`RANDOM}};
  mesh_8_8_io_in_control_0_dataflow_pipe_b = _RAND_2353[0:0];
  _RAND_2354 = {1{`RANDOM}};
  mesh_8_8_io_in_control_0_propagate_pipe_b = _RAND_2354[0:0];
  _RAND_2355 = {1{`RANDOM}};
  mesh_8_8_io_in_control_1_shift_pipe_b = _RAND_2355[4:0];
  _RAND_2356 = {1{`RANDOM}};
  mesh_8_8_io_in_control_1_dataflow_pipe_b = _RAND_2356[0:0];
  _RAND_2357 = {1{`RANDOM}};
  mesh_8_8_io_in_control_1_propagate_pipe_b = _RAND_2357[0:0];
  _RAND_2358 = {1{`RANDOM}};
  mesh_9_8_io_in_control_0_shift_pipe_b = _RAND_2358[4:0];
  _RAND_2359 = {1{`RANDOM}};
  mesh_9_8_io_in_control_0_dataflow_pipe_b = _RAND_2359[0:0];
  _RAND_2360 = {1{`RANDOM}};
  mesh_9_8_io_in_control_0_propagate_pipe_b = _RAND_2360[0:0];
  _RAND_2361 = {1{`RANDOM}};
  mesh_9_8_io_in_control_1_shift_pipe_b = _RAND_2361[4:0];
  _RAND_2362 = {1{`RANDOM}};
  mesh_9_8_io_in_control_1_dataflow_pipe_b = _RAND_2362[0:0];
  _RAND_2363 = {1{`RANDOM}};
  mesh_9_8_io_in_control_1_propagate_pipe_b = _RAND_2363[0:0];
  _RAND_2364 = {1{`RANDOM}};
  mesh_10_8_io_in_control_0_shift_pipe_b = _RAND_2364[4:0];
  _RAND_2365 = {1{`RANDOM}};
  mesh_10_8_io_in_control_0_dataflow_pipe_b = _RAND_2365[0:0];
  _RAND_2366 = {1{`RANDOM}};
  mesh_10_8_io_in_control_0_propagate_pipe_b = _RAND_2366[0:0];
  _RAND_2367 = {1{`RANDOM}};
  mesh_10_8_io_in_control_1_shift_pipe_b = _RAND_2367[4:0];
  _RAND_2368 = {1{`RANDOM}};
  mesh_10_8_io_in_control_1_dataflow_pipe_b = _RAND_2368[0:0];
  _RAND_2369 = {1{`RANDOM}};
  mesh_10_8_io_in_control_1_propagate_pipe_b = _RAND_2369[0:0];
  _RAND_2370 = {1{`RANDOM}};
  mesh_11_8_io_in_control_0_shift_pipe_b = _RAND_2370[4:0];
  _RAND_2371 = {1{`RANDOM}};
  mesh_11_8_io_in_control_0_dataflow_pipe_b = _RAND_2371[0:0];
  _RAND_2372 = {1{`RANDOM}};
  mesh_11_8_io_in_control_0_propagate_pipe_b = _RAND_2372[0:0];
  _RAND_2373 = {1{`RANDOM}};
  mesh_11_8_io_in_control_1_shift_pipe_b = _RAND_2373[4:0];
  _RAND_2374 = {1{`RANDOM}};
  mesh_11_8_io_in_control_1_dataflow_pipe_b = _RAND_2374[0:0];
  _RAND_2375 = {1{`RANDOM}};
  mesh_11_8_io_in_control_1_propagate_pipe_b = _RAND_2375[0:0];
  _RAND_2376 = {1{`RANDOM}};
  mesh_12_8_io_in_control_0_shift_pipe_b = _RAND_2376[4:0];
  _RAND_2377 = {1{`RANDOM}};
  mesh_12_8_io_in_control_0_dataflow_pipe_b = _RAND_2377[0:0];
  _RAND_2378 = {1{`RANDOM}};
  mesh_12_8_io_in_control_0_propagate_pipe_b = _RAND_2378[0:0];
  _RAND_2379 = {1{`RANDOM}};
  mesh_12_8_io_in_control_1_shift_pipe_b = _RAND_2379[4:0];
  _RAND_2380 = {1{`RANDOM}};
  mesh_12_8_io_in_control_1_dataflow_pipe_b = _RAND_2380[0:0];
  _RAND_2381 = {1{`RANDOM}};
  mesh_12_8_io_in_control_1_propagate_pipe_b = _RAND_2381[0:0];
  _RAND_2382 = {1{`RANDOM}};
  mesh_13_8_io_in_control_0_shift_pipe_b = _RAND_2382[4:0];
  _RAND_2383 = {1{`RANDOM}};
  mesh_13_8_io_in_control_0_dataflow_pipe_b = _RAND_2383[0:0];
  _RAND_2384 = {1{`RANDOM}};
  mesh_13_8_io_in_control_0_propagate_pipe_b = _RAND_2384[0:0];
  _RAND_2385 = {1{`RANDOM}};
  mesh_13_8_io_in_control_1_shift_pipe_b = _RAND_2385[4:0];
  _RAND_2386 = {1{`RANDOM}};
  mesh_13_8_io_in_control_1_dataflow_pipe_b = _RAND_2386[0:0];
  _RAND_2387 = {1{`RANDOM}};
  mesh_13_8_io_in_control_1_propagate_pipe_b = _RAND_2387[0:0];
  _RAND_2388 = {1{`RANDOM}};
  mesh_14_8_io_in_control_0_shift_pipe_b = _RAND_2388[4:0];
  _RAND_2389 = {1{`RANDOM}};
  mesh_14_8_io_in_control_0_dataflow_pipe_b = _RAND_2389[0:0];
  _RAND_2390 = {1{`RANDOM}};
  mesh_14_8_io_in_control_0_propagate_pipe_b = _RAND_2390[0:0];
  _RAND_2391 = {1{`RANDOM}};
  mesh_14_8_io_in_control_1_shift_pipe_b = _RAND_2391[4:0];
  _RAND_2392 = {1{`RANDOM}};
  mesh_14_8_io_in_control_1_dataflow_pipe_b = _RAND_2392[0:0];
  _RAND_2393 = {1{`RANDOM}};
  mesh_14_8_io_in_control_1_propagate_pipe_b = _RAND_2393[0:0];
  _RAND_2394 = {1{`RANDOM}};
  mesh_15_8_io_in_control_0_shift_pipe_b = _RAND_2394[4:0];
  _RAND_2395 = {1{`RANDOM}};
  mesh_15_8_io_in_control_0_dataflow_pipe_b = _RAND_2395[0:0];
  _RAND_2396 = {1{`RANDOM}};
  mesh_15_8_io_in_control_0_propagate_pipe_b = _RAND_2396[0:0];
  _RAND_2397 = {1{`RANDOM}};
  mesh_15_8_io_in_control_1_shift_pipe_b = _RAND_2397[4:0];
  _RAND_2398 = {1{`RANDOM}};
  mesh_15_8_io_in_control_1_dataflow_pipe_b = _RAND_2398[0:0];
  _RAND_2399 = {1{`RANDOM}};
  mesh_15_8_io_in_control_1_propagate_pipe_b = _RAND_2399[0:0];
  _RAND_2400 = {1{`RANDOM}};
  mesh_0_9_io_in_control_0_shift_pipe_b = _RAND_2400[4:0];
  _RAND_2401 = {1{`RANDOM}};
  mesh_0_9_io_in_control_0_dataflow_pipe_b = _RAND_2401[0:0];
  _RAND_2402 = {1{`RANDOM}};
  mesh_0_9_io_in_control_0_propagate_pipe_b = _RAND_2402[0:0];
  _RAND_2403 = {1{`RANDOM}};
  mesh_0_9_io_in_control_1_shift_pipe_b = _RAND_2403[4:0];
  _RAND_2404 = {1{`RANDOM}};
  mesh_0_9_io_in_control_1_dataflow_pipe_b = _RAND_2404[0:0];
  _RAND_2405 = {1{`RANDOM}};
  mesh_0_9_io_in_control_1_propagate_pipe_b = _RAND_2405[0:0];
  _RAND_2406 = {1{`RANDOM}};
  mesh_1_9_io_in_control_0_shift_pipe_b = _RAND_2406[4:0];
  _RAND_2407 = {1{`RANDOM}};
  mesh_1_9_io_in_control_0_dataflow_pipe_b = _RAND_2407[0:0];
  _RAND_2408 = {1{`RANDOM}};
  mesh_1_9_io_in_control_0_propagate_pipe_b = _RAND_2408[0:0];
  _RAND_2409 = {1{`RANDOM}};
  mesh_1_9_io_in_control_1_shift_pipe_b = _RAND_2409[4:0];
  _RAND_2410 = {1{`RANDOM}};
  mesh_1_9_io_in_control_1_dataflow_pipe_b = _RAND_2410[0:0];
  _RAND_2411 = {1{`RANDOM}};
  mesh_1_9_io_in_control_1_propagate_pipe_b = _RAND_2411[0:0];
  _RAND_2412 = {1{`RANDOM}};
  mesh_2_9_io_in_control_0_shift_pipe_b = _RAND_2412[4:0];
  _RAND_2413 = {1{`RANDOM}};
  mesh_2_9_io_in_control_0_dataflow_pipe_b = _RAND_2413[0:0];
  _RAND_2414 = {1{`RANDOM}};
  mesh_2_9_io_in_control_0_propagate_pipe_b = _RAND_2414[0:0];
  _RAND_2415 = {1{`RANDOM}};
  mesh_2_9_io_in_control_1_shift_pipe_b = _RAND_2415[4:0];
  _RAND_2416 = {1{`RANDOM}};
  mesh_2_9_io_in_control_1_dataflow_pipe_b = _RAND_2416[0:0];
  _RAND_2417 = {1{`RANDOM}};
  mesh_2_9_io_in_control_1_propagate_pipe_b = _RAND_2417[0:0];
  _RAND_2418 = {1{`RANDOM}};
  mesh_3_9_io_in_control_0_shift_pipe_b = _RAND_2418[4:0];
  _RAND_2419 = {1{`RANDOM}};
  mesh_3_9_io_in_control_0_dataflow_pipe_b = _RAND_2419[0:0];
  _RAND_2420 = {1{`RANDOM}};
  mesh_3_9_io_in_control_0_propagate_pipe_b = _RAND_2420[0:0];
  _RAND_2421 = {1{`RANDOM}};
  mesh_3_9_io_in_control_1_shift_pipe_b = _RAND_2421[4:0];
  _RAND_2422 = {1{`RANDOM}};
  mesh_3_9_io_in_control_1_dataflow_pipe_b = _RAND_2422[0:0];
  _RAND_2423 = {1{`RANDOM}};
  mesh_3_9_io_in_control_1_propagate_pipe_b = _RAND_2423[0:0];
  _RAND_2424 = {1{`RANDOM}};
  mesh_4_9_io_in_control_0_shift_pipe_b = _RAND_2424[4:0];
  _RAND_2425 = {1{`RANDOM}};
  mesh_4_9_io_in_control_0_dataflow_pipe_b = _RAND_2425[0:0];
  _RAND_2426 = {1{`RANDOM}};
  mesh_4_9_io_in_control_0_propagate_pipe_b = _RAND_2426[0:0];
  _RAND_2427 = {1{`RANDOM}};
  mesh_4_9_io_in_control_1_shift_pipe_b = _RAND_2427[4:0];
  _RAND_2428 = {1{`RANDOM}};
  mesh_4_9_io_in_control_1_dataflow_pipe_b = _RAND_2428[0:0];
  _RAND_2429 = {1{`RANDOM}};
  mesh_4_9_io_in_control_1_propagate_pipe_b = _RAND_2429[0:0];
  _RAND_2430 = {1{`RANDOM}};
  mesh_5_9_io_in_control_0_shift_pipe_b = _RAND_2430[4:0];
  _RAND_2431 = {1{`RANDOM}};
  mesh_5_9_io_in_control_0_dataflow_pipe_b = _RAND_2431[0:0];
  _RAND_2432 = {1{`RANDOM}};
  mesh_5_9_io_in_control_0_propagate_pipe_b = _RAND_2432[0:0];
  _RAND_2433 = {1{`RANDOM}};
  mesh_5_9_io_in_control_1_shift_pipe_b = _RAND_2433[4:0];
  _RAND_2434 = {1{`RANDOM}};
  mesh_5_9_io_in_control_1_dataflow_pipe_b = _RAND_2434[0:0];
  _RAND_2435 = {1{`RANDOM}};
  mesh_5_9_io_in_control_1_propagate_pipe_b = _RAND_2435[0:0];
  _RAND_2436 = {1{`RANDOM}};
  mesh_6_9_io_in_control_0_shift_pipe_b = _RAND_2436[4:0];
  _RAND_2437 = {1{`RANDOM}};
  mesh_6_9_io_in_control_0_dataflow_pipe_b = _RAND_2437[0:0];
  _RAND_2438 = {1{`RANDOM}};
  mesh_6_9_io_in_control_0_propagate_pipe_b = _RAND_2438[0:0];
  _RAND_2439 = {1{`RANDOM}};
  mesh_6_9_io_in_control_1_shift_pipe_b = _RAND_2439[4:0];
  _RAND_2440 = {1{`RANDOM}};
  mesh_6_9_io_in_control_1_dataflow_pipe_b = _RAND_2440[0:0];
  _RAND_2441 = {1{`RANDOM}};
  mesh_6_9_io_in_control_1_propagate_pipe_b = _RAND_2441[0:0];
  _RAND_2442 = {1{`RANDOM}};
  mesh_7_9_io_in_control_0_shift_pipe_b = _RAND_2442[4:0];
  _RAND_2443 = {1{`RANDOM}};
  mesh_7_9_io_in_control_0_dataflow_pipe_b = _RAND_2443[0:0];
  _RAND_2444 = {1{`RANDOM}};
  mesh_7_9_io_in_control_0_propagate_pipe_b = _RAND_2444[0:0];
  _RAND_2445 = {1{`RANDOM}};
  mesh_7_9_io_in_control_1_shift_pipe_b = _RAND_2445[4:0];
  _RAND_2446 = {1{`RANDOM}};
  mesh_7_9_io_in_control_1_dataflow_pipe_b = _RAND_2446[0:0];
  _RAND_2447 = {1{`RANDOM}};
  mesh_7_9_io_in_control_1_propagate_pipe_b = _RAND_2447[0:0];
  _RAND_2448 = {1{`RANDOM}};
  mesh_8_9_io_in_control_0_shift_pipe_b = _RAND_2448[4:0];
  _RAND_2449 = {1{`RANDOM}};
  mesh_8_9_io_in_control_0_dataflow_pipe_b = _RAND_2449[0:0];
  _RAND_2450 = {1{`RANDOM}};
  mesh_8_9_io_in_control_0_propagate_pipe_b = _RAND_2450[0:0];
  _RAND_2451 = {1{`RANDOM}};
  mesh_8_9_io_in_control_1_shift_pipe_b = _RAND_2451[4:0];
  _RAND_2452 = {1{`RANDOM}};
  mesh_8_9_io_in_control_1_dataflow_pipe_b = _RAND_2452[0:0];
  _RAND_2453 = {1{`RANDOM}};
  mesh_8_9_io_in_control_1_propagate_pipe_b = _RAND_2453[0:0];
  _RAND_2454 = {1{`RANDOM}};
  mesh_9_9_io_in_control_0_shift_pipe_b = _RAND_2454[4:0];
  _RAND_2455 = {1{`RANDOM}};
  mesh_9_9_io_in_control_0_dataflow_pipe_b = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  mesh_9_9_io_in_control_0_propagate_pipe_b = _RAND_2456[0:0];
  _RAND_2457 = {1{`RANDOM}};
  mesh_9_9_io_in_control_1_shift_pipe_b = _RAND_2457[4:0];
  _RAND_2458 = {1{`RANDOM}};
  mesh_9_9_io_in_control_1_dataflow_pipe_b = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  mesh_9_9_io_in_control_1_propagate_pipe_b = _RAND_2459[0:0];
  _RAND_2460 = {1{`RANDOM}};
  mesh_10_9_io_in_control_0_shift_pipe_b = _RAND_2460[4:0];
  _RAND_2461 = {1{`RANDOM}};
  mesh_10_9_io_in_control_0_dataflow_pipe_b = _RAND_2461[0:0];
  _RAND_2462 = {1{`RANDOM}};
  mesh_10_9_io_in_control_0_propagate_pipe_b = _RAND_2462[0:0];
  _RAND_2463 = {1{`RANDOM}};
  mesh_10_9_io_in_control_1_shift_pipe_b = _RAND_2463[4:0];
  _RAND_2464 = {1{`RANDOM}};
  mesh_10_9_io_in_control_1_dataflow_pipe_b = _RAND_2464[0:0];
  _RAND_2465 = {1{`RANDOM}};
  mesh_10_9_io_in_control_1_propagate_pipe_b = _RAND_2465[0:0];
  _RAND_2466 = {1{`RANDOM}};
  mesh_11_9_io_in_control_0_shift_pipe_b = _RAND_2466[4:0];
  _RAND_2467 = {1{`RANDOM}};
  mesh_11_9_io_in_control_0_dataflow_pipe_b = _RAND_2467[0:0];
  _RAND_2468 = {1{`RANDOM}};
  mesh_11_9_io_in_control_0_propagate_pipe_b = _RAND_2468[0:0];
  _RAND_2469 = {1{`RANDOM}};
  mesh_11_9_io_in_control_1_shift_pipe_b = _RAND_2469[4:0];
  _RAND_2470 = {1{`RANDOM}};
  mesh_11_9_io_in_control_1_dataflow_pipe_b = _RAND_2470[0:0];
  _RAND_2471 = {1{`RANDOM}};
  mesh_11_9_io_in_control_1_propagate_pipe_b = _RAND_2471[0:0];
  _RAND_2472 = {1{`RANDOM}};
  mesh_12_9_io_in_control_0_shift_pipe_b = _RAND_2472[4:0];
  _RAND_2473 = {1{`RANDOM}};
  mesh_12_9_io_in_control_0_dataflow_pipe_b = _RAND_2473[0:0];
  _RAND_2474 = {1{`RANDOM}};
  mesh_12_9_io_in_control_0_propagate_pipe_b = _RAND_2474[0:0];
  _RAND_2475 = {1{`RANDOM}};
  mesh_12_9_io_in_control_1_shift_pipe_b = _RAND_2475[4:0];
  _RAND_2476 = {1{`RANDOM}};
  mesh_12_9_io_in_control_1_dataflow_pipe_b = _RAND_2476[0:0];
  _RAND_2477 = {1{`RANDOM}};
  mesh_12_9_io_in_control_1_propagate_pipe_b = _RAND_2477[0:0];
  _RAND_2478 = {1{`RANDOM}};
  mesh_13_9_io_in_control_0_shift_pipe_b = _RAND_2478[4:0];
  _RAND_2479 = {1{`RANDOM}};
  mesh_13_9_io_in_control_0_dataflow_pipe_b = _RAND_2479[0:0];
  _RAND_2480 = {1{`RANDOM}};
  mesh_13_9_io_in_control_0_propagate_pipe_b = _RAND_2480[0:0];
  _RAND_2481 = {1{`RANDOM}};
  mesh_13_9_io_in_control_1_shift_pipe_b = _RAND_2481[4:0];
  _RAND_2482 = {1{`RANDOM}};
  mesh_13_9_io_in_control_1_dataflow_pipe_b = _RAND_2482[0:0];
  _RAND_2483 = {1{`RANDOM}};
  mesh_13_9_io_in_control_1_propagate_pipe_b = _RAND_2483[0:0];
  _RAND_2484 = {1{`RANDOM}};
  mesh_14_9_io_in_control_0_shift_pipe_b = _RAND_2484[4:0];
  _RAND_2485 = {1{`RANDOM}};
  mesh_14_9_io_in_control_0_dataflow_pipe_b = _RAND_2485[0:0];
  _RAND_2486 = {1{`RANDOM}};
  mesh_14_9_io_in_control_0_propagate_pipe_b = _RAND_2486[0:0];
  _RAND_2487 = {1{`RANDOM}};
  mesh_14_9_io_in_control_1_shift_pipe_b = _RAND_2487[4:0];
  _RAND_2488 = {1{`RANDOM}};
  mesh_14_9_io_in_control_1_dataflow_pipe_b = _RAND_2488[0:0];
  _RAND_2489 = {1{`RANDOM}};
  mesh_14_9_io_in_control_1_propagate_pipe_b = _RAND_2489[0:0];
  _RAND_2490 = {1{`RANDOM}};
  mesh_15_9_io_in_control_0_shift_pipe_b = _RAND_2490[4:0];
  _RAND_2491 = {1{`RANDOM}};
  mesh_15_9_io_in_control_0_dataflow_pipe_b = _RAND_2491[0:0];
  _RAND_2492 = {1{`RANDOM}};
  mesh_15_9_io_in_control_0_propagate_pipe_b = _RAND_2492[0:0];
  _RAND_2493 = {1{`RANDOM}};
  mesh_15_9_io_in_control_1_shift_pipe_b = _RAND_2493[4:0];
  _RAND_2494 = {1{`RANDOM}};
  mesh_15_9_io_in_control_1_dataflow_pipe_b = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  mesh_15_9_io_in_control_1_propagate_pipe_b = _RAND_2495[0:0];
  _RAND_2496 = {1{`RANDOM}};
  mesh_0_10_io_in_control_0_shift_pipe_b = _RAND_2496[4:0];
  _RAND_2497 = {1{`RANDOM}};
  mesh_0_10_io_in_control_0_dataflow_pipe_b = _RAND_2497[0:0];
  _RAND_2498 = {1{`RANDOM}};
  mesh_0_10_io_in_control_0_propagate_pipe_b = _RAND_2498[0:0];
  _RAND_2499 = {1{`RANDOM}};
  mesh_0_10_io_in_control_1_shift_pipe_b = _RAND_2499[4:0];
  _RAND_2500 = {1{`RANDOM}};
  mesh_0_10_io_in_control_1_dataflow_pipe_b = _RAND_2500[0:0];
  _RAND_2501 = {1{`RANDOM}};
  mesh_0_10_io_in_control_1_propagate_pipe_b = _RAND_2501[0:0];
  _RAND_2502 = {1{`RANDOM}};
  mesh_1_10_io_in_control_0_shift_pipe_b = _RAND_2502[4:0];
  _RAND_2503 = {1{`RANDOM}};
  mesh_1_10_io_in_control_0_dataflow_pipe_b = _RAND_2503[0:0];
  _RAND_2504 = {1{`RANDOM}};
  mesh_1_10_io_in_control_0_propagate_pipe_b = _RAND_2504[0:0];
  _RAND_2505 = {1{`RANDOM}};
  mesh_1_10_io_in_control_1_shift_pipe_b = _RAND_2505[4:0];
  _RAND_2506 = {1{`RANDOM}};
  mesh_1_10_io_in_control_1_dataflow_pipe_b = _RAND_2506[0:0];
  _RAND_2507 = {1{`RANDOM}};
  mesh_1_10_io_in_control_1_propagate_pipe_b = _RAND_2507[0:0];
  _RAND_2508 = {1{`RANDOM}};
  mesh_2_10_io_in_control_0_shift_pipe_b = _RAND_2508[4:0];
  _RAND_2509 = {1{`RANDOM}};
  mesh_2_10_io_in_control_0_dataflow_pipe_b = _RAND_2509[0:0];
  _RAND_2510 = {1{`RANDOM}};
  mesh_2_10_io_in_control_0_propagate_pipe_b = _RAND_2510[0:0];
  _RAND_2511 = {1{`RANDOM}};
  mesh_2_10_io_in_control_1_shift_pipe_b = _RAND_2511[4:0];
  _RAND_2512 = {1{`RANDOM}};
  mesh_2_10_io_in_control_1_dataflow_pipe_b = _RAND_2512[0:0];
  _RAND_2513 = {1{`RANDOM}};
  mesh_2_10_io_in_control_1_propagate_pipe_b = _RAND_2513[0:0];
  _RAND_2514 = {1{`RANDOM}};
  mesh_3_10_io_in_control_0_shift_pipe_b = _RAND_2514[4:0];
  _RAND_2515 = {1{`RANDOM}};
  mesh_3_10_io_in_control_0_dataflow_pipe_b = _RAND_2515[0:0];
  _RAND_2516 = {1{`RANDOM}};
  mesh_3_10_io_in_control_0_propagate_pipe_b = _RAND_2516[0:0];
  _RAND_2517 = {1{`RANDOM}};
  mesh_3_10_io_in_control_1_shift_pipe_b = _RAND_2517[4:0];
  _RAND_2518 = {1{`RANDOM}};
  mesh_3_10_io_in_control_1_dataflow_pipe_b = _RAND_2518[0:0];
  _RAND_2519 = {1{`RANDOM}};
  mesh_3_10_io_in_control_1_propagate_pipe_b = _RAND_2519[0:0];
  _RAND_2520 = {1{`RANDOM}};
  mesh_4_10_io_in_control_0_shift_pipe_b = _RAND_2520[4:0];
  _RAND_2521 = {1{`RANDOM}};
  mesh_4_10_io_in_control_0_dataflow_pipe_b = _RAND_2521[0:0];
  _RAND_2522 = {1{`RANDOM}};
  mesh_4_10_io_in_control_0_propagate_pipe_b = _RAND_2522[0:0];
  _RAND_2523 = {1{`RANDOM}};
  mesh_4_10_io_in_control_1_shift_pipe_b = _RAND_2523[4:0];
  _RAND_2524 = {1{`RANDOM}};
  mesh_4_10_io_in_control_1_dataflow_pipe_b = _RAND_2524[0:0];
  _RAND_2525 = {1{`RANDOM}};
  mesh_4_10_io_in_control_1_propagate_pipe_b = _RAND_2525[0:0];
  _RAND_2526 = {1{`RANDOM}};
  mesh_5_10_io_in_control_0_shift_pipe_b = _RAND_2526[4:0];
  _RAND_2527 = {1{`RANDOM}};
  mesh_5_10_io_in_control_0_dataflow_pipe_b = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  mesh_5_10_io_in_control_0_propagate_pipe_b = _RAND_2528[0:0];
  _RAND_2529 = {1{`RANDOM}};
  mesh_5_10_io_in_control_1_shift_pipe_b = _RAND_2529[4:0];
  _RAND_2530 = {1{`RANDOM}};
  mesh_5_10_io_in_control_1_dataflow_pipe_b = _RAND_2530[0:0];
  _RAND_2531 = {1{`RANDOM}};
  mesh_5_10_io_in_control_1_propagate_pipe_b = _RAND_2531[0:0];
  _RAND_2532 = {1{`RANDOM}};
  mesh_6_10_io_in_control_0_shift_pipe_b = _RAND_2532[4:0];
  _RAND_2533 = {1{`RANDOM}};
  mesh_6_10_io_in_control_0_dataflow_pipe_b = _RAND_2533[0:0];
  _RAND_2534 = {1{`RANDOM}};
  mesh_6_10_io_in_control_0_propagate_pipe_b = _RAND_2534[0:0];
  _RAND_2535 = {1{`RANDOM}};
  mesh_6_10_io_in_control_1_shift_pipe_b = _RAND_2535[4:0];
  _RAND_2536 = {1{`RANDOM}};
  mesh_6_10_io_in_control_1_dataflow_pipe_b = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  mesh_6_10_io_in_control_1_propagate_pipe_b = _RAND_2537[0:0];
  _RAND_2538 = {1{`RANDOM}};
  mesh_7_10_io_in_control_0_shift_pipe_b = _RAND_2538[4:0];
  _RAND_2539 = {1{`RANDOM}};
  mesh_7_10_io_in_control_0_dataflow_pipe_b = _RAND_2539[0:0];
  _RAND_2540 = {1{`RANDOM}};
  mesh_7_10_io_in_control_0_propagate_pipe_b = _RAND_2540[0:0];
  _RAND_2541 = {1{`RANDOM}};
  mesh_7_10_io_in_control_1_shift_pipe_b = _RAND_2541[4:0];
  _RAND_2542 = {1{`RANDOM}};
  mesh_7_10_io_in_control_1_dataflow_pipe_b = _RAND_2542[0:0];
  _RAND_2543 = {1{`RANDOM}};
  mesh_7_10_io_in_control_1_propagate_pipe_b = _RAND_2543[0:0];
  _RAND_2544 = {1{`RANDOM}};
  mesh_8_10_io_in_control_0_shift_pipe_b = _RAND_2544[4:0];
  _RAND_2545 = {1{`RANDOM}};
  mesh_8_10_io_in_control_0_dataflow_pipe_b = _RAND_2545[0:0];
  _RAND_2546 = {1{`RANDOM}};
  mesh_8_10_io_in_control_0_propagate_pipe_b = _RAND_2546[0:0];
  _RAND_2547 = {1{`RANDOM}};
  mesh_8_10_io_in_control_1_shift_pipe_b = _RAND_2547[4:0];
  _RAND_2548 = {1{`RANDOM}};
  mesh_8_10_io_in_control_1_dataflow_pipe_b = _RAND_2548[0:0];
  _RAND_2549 = {1{`RANDOM}};
  mesh_8_10_io_in_control_1_propagate_pipe_b = _RAND_2549[0:0];
  _RAND_2550 = {1{`RANDOM}};
  mesh_9_10_io_in_control_0_shift_pipe_b = _RAND_2550[4:0];
  _RAND_2551 = {1{`RANDOM}};
  mesh_9_10_io_in_control_0_dataflow_pipe_b = _RAND_2551[0:0];
  _RAND_2552 = {1{`RANDOM}};
  mesh_9_10_io_in_control_0_propagate_pipe_b = _RAND_2552[0:0];
  _RAND_2553 = {1{`RANDOM}};
  mesh_9_10_io_in_control_1_shift_pipe_b = _RAND_2553[4:0];
  _RAND_2554 = {1{`RANDOM}};
  mesh_9_10_io_in_control_1_dataflow_pipe_b = _RAND_2554[0:0];
  _RAND_2555 = {1{`RANDOM}};
  mesh_9_10_io_in_control_1_propagate_pipe_b = _RAND_2555[0:0];
  _RAND_2556 = {1{`RANDOM}};
  mesh_10_10_io_in_control_0_shift_pipe_b = _RAND_2556[4:0];
  _RAND_2557 = {1{`RANDOM}};
  mesh_10_10_io_in_control_0_dataflow_pipe_b = _RAND_2557[0:0];
  _RAND_2558 = {1{`RANDOM}};
  mesh_10_10_io_in_control_0_propagate_pipe_b = _RAND_2558[0:0];
  _RAND_2559 = {1{`RANDOM}};
  mesh_10_10_io_in_control_1_shift_pipe_b = _RAND_2559[4:0];
  _RAND_2560 = {1{`RANDOM}};
  mesh_10_10_io_in_control_1_dataflow_pipe_b = _RAND_2560[0:0];
  _RAND_2561 = {1{`RANDOM}};
  mesh_10_10_io_in_control_1_propagate_pipe_b = _RAND_2561[0:0];
  _RAND_2562 = {1{`RANDOM}};
  mesh_11_10_io_in_control_0_shift_pipe_b = _RAND_2562[4:0];
  _RAND_2563 = {1{`RANDOM}};
  mesh_11_10_io_in_control_0_dataflow_pipe_b = _RAND_2563[0:0];
  _RAND_2564 = {1{`RANDOM}};
  mesh_11_10_io_in_control_0_propagate_pipe_b = _RAND_2564[0:0];
  _RAND_2565 = {1{`RANDOM}};
  mesh_11_10_io_in_control_1_shift_pipe_b = _RAND_2565[4:0];
  _RAND_2566 = {1{`RANDOM}};
  mesh_11_10_io_in_control_1_dataflow_pipe_b = _RAND_2566[0:0];
  _RAND_2567 = {1{`RANDOM}};
  mesh_11_10_io_in_control_1_propagate_pipe_b = _RAND_2567[0:0];
  _RAND_2568 = {1{`RANDOM}};
  mesh_12_10_io_in_control_0_shift_pipe_b = _RAND_2568[4:0];
  _RAND_2569 = {1{`RANDOM}};
  mesh_12_10_io_in_control_0_dataflow_pipe_b = _RAND_2569[0:0];
  _RAND_2570 = {1{`RANDOM}};
  mesh_12_10_io_in_control_0_propagate_pipe_b = _RAND_2570[0:0];
  _RAND_2571 = {1{`RANDOM}};
  mesh_12_10_io_in_control_1_shift_pipe_b = _RAND_2571[4:0];
  _RAND_2572 = {1{`RANDOM}};
  mesh_12_10_io_in_control_1_dataflow_pipe_b = _RAND_2572[0:0];
  _RAND_2573 = {1{`RANDOM}};
  mesh_12_10_io_in_control_1_propagate_pipe_b = _RAND_2573[0:0];
  _RAND_2574 = {1{`RANDOM}};
  mesh_13_10_io_in_control_0_shift_pipe_b = _RAND_2574[4:0];
  _RAND_2575 = {1{`RANDOM}};
  mesh_13_10_io_in_control_0_dataflow_pipe_b = _RAND_2575[0:0];
  _RAND_2576 = {1{`RANDOM}};
  mesh_13_10_io_in_control_0_propagate_pipe_b = _RAND_2576[0:0];
  _RAND_2577 = {1{`RANDOM}};
  mesh_13_10_io_in_control_1_shift_pipe_b = _RAND_2577[4:0];
  _RAND_2578 = {1{`RANDOM}};
  mesh_13_10_io_in_control_1_dataflow_pipe_b = _RAND_2578[0:0];
  _RAND_2579 = {1{`RANDOM}};
  mesh_13_10_io_in_control_1_propagate_pipe_b = _RAND_2579[0:0];
  _RAND_2580 = {1{`RANDOM}};
  mesh_14_10_io_in_control_0_shift_pipe_b = _RAND_2580[4:0];
  _RAND_2581 = {1{`RANDOM}};
  mesh_14_10_io_in_control_0_dataflow_pipe_b = _RAND_2581[0:0];
  _RAND_2582 = {1{`RANDOM}};
  mesh_14_10_io_in_control_0_propagate_pipe_b = _RAND_2582[0:0];
  _RAND_2583 = {1{`RANDOM}};
  mesh_14_10_io_in_control_1_shift_pipe_b = _RAND_2583[4:0];
  _RAND_2584 = {1{`RANDOM}};
  mesh_14_10_io_in_control_1_dataflow_pipe_b = _RAND_2584[0:0];
  _RAND_2585 = {1{`RANDOM}};
  mesh_14_10_io_in_control_1_propagate_pipe_b = _RAND_2585[0:0];
  _RAND_2586 = {1{`RANDOM}};
  mesh_15_10_io_in_control_0_shift_pipe_b = _RAND_2586[4:0];
  _RAND_2587 = {1{`RANDOM}};
  mesh_15_10_io_in_control_0_dataflow_pipe_b = _RAND_2587[0:0];
  _RAND_2588 = {1{`RANDOM}};
  mesh_15_10_io_in_control_0_propagate_pipe_b = _RAND_2588[0:0];
  _RAND_2589 = {1{`RANDOM}};
  mesh_15_10_io_in_control_1_shift_pipe_b = _RAND_2589[4:0];
  _RAND_2590 = {1{`RANDOM}};
  mesh_15_10_io_in_control_1_dataflow_pipe_b = _RAND_2590[0:0];
  _RAND_2591 = {1{`RANDOM}};
  mesh_15_10_io_in_control_1_propagate_pipe_b = _RAND_2591[0:0];
  _RAND_2592 = {1{`RANDOM}};
  mesh_0_11_io_in_control_0_shift_pipe_b = _RAND_2592[4:0];
  _RAND_2593 = {1{`RANDOM}};
  mesh_0_11_io_in_control_0_dataflow_pipe_b = _RAND_2593[0:0];
  _RAND_2594 = {1{`RANDOM}};
  mesh_0_11_io_in_control_0_propagate_pipe_b = _RAND_2594[0:0];
  _RAND_2595 = {1{`RANDOM}};
  mesh_0_11_io_in_control_1_shift_pipe_b = _RAND_2595[4:0];
  _RAND_2596 = {1{`RANDOM}};
  mesh_0_11_io_in_control_1_dataflow_pipe_b = _RAND_2596[0:0];
  _RAND_2597 = {1{`RANDOM}};
  mesh_0_11_io_in_control_1_propagate_pipe_b = _RAND_2597[0:0];
  _RAND_2598 = {1{`RANDOM}};
  mesh_1_11_io_in_control_0_shift_pipe_b = _RAND_2598[4:0];
  _RAND_2599 = {1{`RANDOM}};
  mesh_1_11_io_in_control_0_dataflow_pipe_b = _RAND_2599[0:0];
  _RAND_2600 = {1{`RANDOM}};
  mesh_1_11_io_in_control_0_propagate_pipe_b = _RAND_2600[0:0];
  _RAND_2601 = {1{`RANDOM}};
  mesh_1_11_io_in_control_1_shift_pipe_b = _RAND_2601[4:0];
  _RAND_2602 = {1{`RANDOM}};
  mesh_1_11_io_in_control_1_dataflow_pipe_b = _RAND_2602[0:0];
  _RAND_2603 = {1{`RANDOM}};
  mesh_1_11_io_in_control_1_propagate_pipe_b = _RAND_2603[0:0];
  _RAND_2604 = {1{`RANDOM}};
  mesh_2_11_io_in_control_0_shift_pipe_b = _RAND_2604[4:0];
  _RAND_2605 = {1{`RANDOM}};
  mesh_2_11_io_in_control_0_dataflow_pipe_b = _RAND_2605[0:0];
  _RAND_2606 = {1{`RANDOM}};
  mesh_2_11_io_in_control_0_propagate_pipe_b = _RAND_2606[0:0];
  _RAND_2607 = {1{`RANDOM}};
  mesh_2_11_io_in_control_1_shift_pipe_b = _RAND_2607[4:0];
  _RAND_2608 = {1{`RANDOM}};
  mesh_2_11_io_in_control_1_dataflow_pipe_b = _RAND_2608[0:0];
  _RAND_2609 = {1{`RANDOM}};
  mesh_2_11_io_in_control_1_propagate_pipe_b = _RAND_2609[0:0];
  _RAND_2610 = {1{`RANDOM}};
  mesh_3_11_io_in_control_0_shift_pipe_b = _RAND_2610[4:0];
  _RAND_2611 = {1{`RANDOM}};
  mesh_3_11_io_in_control_0_dataflow_pipe_b = _RAND_2611[0:0];
  _RAND_2612 = {1{`RANDOM}};
  mesh_3_11_io_in_control_0_propagate_pipe_b = _RAND_2612[0:0];
  _RAND_2613 = {1{`RANDOM}};
  mesh_3_11_io_in_control_1_shift_pipe_b = _RAND_2613[4:0];
  _RAND_2614 = {1{`RANDOM}};
  mesh_3_11_io_in_control_1_dataflow_pipe_b = _RAND_2614[0:0];
  _RAND_2615 = {1{`RANDOM}};
  mesh_3_11_io_in_control_1_propagate_pipe_b = _RAND_2615[0:0];
  _RAND_2616 = {1{`RANDOM}};
  mesh_4_11_io_in_control_0_shift_pipe_b = _RAND_2616[4:0];
  _RAND_2617 = {1{`RANDOM}};
  mesh_4_11_io_in_control_0_dataflow_pipe_b = _RAND_2617[0:0];
  _RAND_2618 = {1{`RANDOM}};
  mesh_4_11_io_in_control_0_propagate_pipe_b = _RAND_2618[0:0];
  _RAND_2619 = {1{`RANDOM}};
  mesh_4_11_io_in_control_1_shift_pipe_b = _RAND_2619[4:0];
  _RAND_2620 = {1{`RANDOM}};
  mesh_4_11_io_in_control_1_dataflow_pipe_b = _RAND_2620[0:0];
  _RAND_2621 = {1{`RANDOM}};
  mesh_4_11_io_in_control_1_propagate_pipe_b = _RAND_2621[0:0];
  _RAND_2622 = {1{`RANDOM}};
  mesh_5_11_io_in_control_0_shift_pipe_b = _RAND_2622[4:0];
  _RAND_2623 = {1{`RANDOM}};
  mesh_5_11_io_in_control_0_dataflow_pipe_b = _RAND_2623[0:0];
  _RAND_2624 = {1{`RANDOM}};
  mesh_5_11_io_in_control_0_propagate_pipe_b = _RAND_2624[0:0];
  _RAND_2625 = {1{`RANDOM}};
  mesh_5_11_io_in_control_1_shift_pipe_b = _RAND_2625[4:0];
  _RAND_2626 = {1{`RANDOM}};
  mesh_5_11_io_in_control_1_dataflow_pipe_b = _RAND_2626[0:0];
  _RAND_2627 = {1{`RANDOM}};
  mesh_5_11_io_in_control_1_propagate_pipe_b = _RAND_2627[0:0];
  _RAND_2628 = {1{`RANDOM}};
  mesh_6_11_io_in_control_0_shift_pipe_b = _RAND_2628[4:0];
  _RAND_2629 = {1{`RANDOM}};
  mesh_6_11_io_in_control_0_dataflow_pipe_b = _RAND_2629[0:0];
  _RAND_2630 = {1{`RANDOM}};
  mesh_6_11_io_in_control_0_propagate_pipe_b = _RAND_2630[0:0];
  _RAND_2631 = {1{`RANDOM}};
  mesh_6_11_io_in_control_1_shift_pipe_b = _RAND_2631[4:0];
  _RAND_2632 = {1{`RANDOM}};
  mesh_6_11_io_in_control_1_dataflow_pipe_b = _RAND_2632[0:0];
  _RAND_2633 = {1{`RANDOM}};
  mesh_6_11_io_in_control_1_propagate_pipe_b = _RAND_2633[0:0];
  _RAND_2634 = {1{`RANDOM}};
  mesh_7_11_io_in_control_0_shift_pipe_b = _RAND_2634[4:0];
  _RAND_2635 = {1{`RANDOM}};
  mesh_7_11_io_in_control_0_dataflow_pipe_b = _RAND_2635[0:0];
  _RAND_2636 = {1{`RANDOM}};
  mesh_7_11_io_in_control_0_propagate_pipe_b = _RAND_2636[0:0];
  _RAND_2637 = {1{`RANDOM}};
  mesh_7_11_io_in_control_1_shift_pipe_b = _RAND_2637[4:0];
  _RAND_2638 = {1{`RANDOM}};
  mesh_7_11_io_in_control_1_dataflow_pipe_b = _RAND_2638[0:0];
  _RAND_2639 = {1{`RANDOM}};
  mesh_7_11_io_in_control_1_propagate_pipe_b = _RAND_2639[0:0];
  _RAND_2640 = {1{`RANDOM}};
  mesh_8_11_io_in_control_0_shift_pipe_b = _RAND_2640[4:0];
  _RAND_2641 = {1{`RANDOM}};
  mesh_8_11_io_in_control_0_dataflow_pipe_b = _RAND_2641[0:0];
  _RAND_2642 = {1{`RANDOM}};
  mesh_8_11_io_in_control_0_propagate_pipe_b = _RAND_2642[0:0];
  _RAND_2643 = {1{`RANDOM}};
  mesh_8_11_io_in_control_1_shift_pipe_b = _RAND_2643[4:0];
  _RAND_2644 = {1{`RANDOM}};
  mesh_8_11_io_in_control_1_dataflow_pipe_b = _RAND_2644[0:0];
  _RAND_2645 = {1{`RANDOM}};
  mesh_8_11_io_in_control_1_propagate_pipe_b = _RAND_2645[0:0];
  _RAND_2646 = {1{`RANDOM}};
  mesh_9_11_io_in_control_0_shift_pipe_b = _RAND_2646[4:0];
  _RAND_2647 = {1{`RANDOM}};
  mesh_9_11_io_in_control_0_dataflow_pipe_b = _RAND_2647[0:0];
  _RAND_2648 = {1{`RANDOM}};
  mesh_9_11_io_in_control_0_propagate_pipe_b = _RAND_2648[0:0];
  _RAND_2649 = {1{`RANDOM}};
  mesh_9_11_io_in_control_1_shift_pipe_b = _RAND_2649[4:0];
  _RAND_2650 = {1{`RANDOM}};
  mesh_9_11_io_in_control_1_dataflow_pipe_b = _RAND_2650[0:0];
  _RAND_2651 = {1{`RANDOM}};
  mesh_9_11_io_in_control_1_propagate_pipe_b = _RAND_2651[0:0];
  _RAND_2652 = {1{`RANDOM}};
  mesh_10_11_io_in_control_0_shift_pipe_b = _RAND_2652[4:0];
  _RAND_2653 = {1{`RANDOM}};
  mesh_10_11_io_in_control_0_dataflow_pipe_b = _RAND_2653[0:0];
  _RAND_2654 = {1{`RANDOM}};
  mesh_10_11_io_in_control_0_propagate_pipe_b = _RAND_2654[0:0];
  _RAND_2655 = {1{`RANDOM}};
  mesh_10_11_io_in_control_1_shift_pipe_b = _RAND_2655[4:0];
  _RAND_2656 = {1{`RANDOM}};
  mesh_10_11_io_in_control_1_dataflow_pipe_b = _RAND_2656[0:0];
  _RAND_2657 = {1{`RANDOM}};
  mesh_10_11_io_in_control_1_propagate_pipe_b = _RAND_2657[0:0];
  _RAND_2658 = {1{`RANDOM}};
  mesh_11_11_io_in_control_0_shift_pipe_b = _RAND_2658[4:0];
  _RAND_2659 = {1{`RANDOM}};
  mesh_11_11_io_in_control_0_dataflow_pipe_b = _RAND_2659[0:0];
  _RAND_2660 = {1{`RANDOM}};
  mesh_11_11_io_in_control_0_propagate_pipe_b = _RAND_2660[0:0];
  _RAND_2661 = {1{`RANDOM}};
  mesh_11_11_io_in_control_1_shift_pipe_b = _RAND_2661[4:0];
  _RAND_2662 = {1{`RANDOM}};
  mesh_11_11_io_in_control_1_dataflow_pipe_b = _RAND_2662[0:0];
  _RAND_2663 = {1{`RANDOM}};
  mesh_11_11_io_in_control_1_propagate_pipe_b = _RAND_2663[0:0];
  _RAND_2664 = {1{`RANDOM}};
  mesh_12_11_io_in_control_0_shift_pipe_b = _RAND_2664[4:0];
  _RAND_2665 = {1{`RANDOM}};
  mesh_12_11_io_in_control_0_dataflow_pipe_b = _RAND_2665[0:0];
  _RAND_2666 = {1{`RANDOM}};
  mesh_12_11_io_in_control_0_propagate_pipe_b = _RAND_2666[0:0];
  _RAND_2667 = {1{`RANDOM}};
  mesh_12_11_io_in_control_1_shift_pipe_b = _RAND_2667[4:0];
  _RAND_2668 = {1{`RANDOM}};
  mesh_12_11_io_in_control_1_dataflow_pipe_b = _RAND_2668[0:0];
  _RAND_2669 = {1{`RANDOM}};
  mesh_12_11_io_in_control_1_propagate_pipe_b = _RAND_2669[0:0];
  _RAND_2670 = {1{`RANDOM}};
  mesh_13_11_io_in_control_0_shift_pipe_b = _RAND_2670[4:0];
  _RAND_2671 = {1{`RANDOM}};
  mesh_13_11_io_in_control_0_dataflow_pipe_b = _RAND_2671[0:0];
  _RAND_2672 = {1{`RANDOM}};
  mesh_13_11_io_in_control_0_propagate_pipe_b = _RAND_2672[0:0];
  _RAND_2673 = {1{`RANDOM}};
  mesh_13_11_io_in_control_1_shift_pipe_b = _RAND_2673[4:0];
  _RAND_2674 = {1{`RANDOM}};
  mesh_13_11_io_in_control_1_dataflow_pipe_b = _RAND_2674[0:0];
  _RAND_2675 = {1{`RANDOM}};
  mesh_13_11_io_in_control_1_propagate_pipe_b = _RAND_2675[0:0];
  _RAND_2676 = {1{`RANDOM}};
  mesh_14_11_io_in_control_0_shift_pipe_b = _RAND_2676[4:0];
  _RAND_2677 = {1{`RANDOM}};
  mesh_14_11_io_in_control_0_dataflow_pipe_b = _RAND_2677[0:0];
  _RAND_2678 = {1{`RANDOM}};
  mesh_14_11_io_in_control_0_propagate_pipe_b = _RAND_2678[0:0];
  _RAND_2679 = {1{`RANDOM}};
  mesh_14_11_io_in_control_1_shift_pipe_b = _RAND_2679[4:0];
  _RAND_2680 = {1{`RANDOM}};
  mesh_14_11_io_in_control_1_dataflow_pipe_b = _RAND_2680[0:0];
  _RAND_2681 = {1{`RANDOM}};
  mesh_14_11_io_in_control_1_propagate_pipe_b = _RAND_2681[0:0];
  _RAND_2682 = {1{`RANDOM}};
  mesh_15_11_io_in_control_0_shift_pipe_b = _RAND_2682[4:0];
  _RAND_2683 = {1{`RANDOM}};
  mesh_15_11_io_in_control_0_dataflow_pipe_b = _RAND_2683[0:0];
  _RAND_2684 = {1{`RANDOM}};
  mesh_15_11_io_in_control_0_propagate_pipe_b = _RAND_2684[0:0];
  _RAND_2685 = {1{`RANDOM}};
  mesh_15_11_io_in_control_1_shift_pipe_b = _RAND_2685[4:0];
  _RAND_2686 = {1{`RANDOM}};
  mesh_15_11_io_in_control_1_dataflow_pipe_b = _RAND_2686[0:0];
  _RAND_2687 = {1{`RANDOM}};
  mesh_15_11_io_in_control_1_propagate_pipe_b = _RAND_2687[0:0];
  _RAND_2688 = {1{`RANDOM}};
  mesh_0_12_io_in_control_0_shift_pipe_b = _RAND_2688[4:0];
  _RAND_2689 = {1{`RANDOM}};
  mesh_0_12_io_in_control_0_dataflow_pipe_b = _RAND_2689[0:0];
  _RAND_2690 = {1{`RANDOM}};
  mesh_0_12_io_in_control_0_propagate_pipe_b = _RAND_2690[0:0];
  _RAND_2691 = {1{`RANDOM}};
  mesh_0_12_io_in_control_1_shift_pipe_b = _RAND_2691[4:0];
  _RAND_2692 = {1{`RANDOM}};
  mesh_0_12_io_in_control_1_dataflow_pipe_b = _RAND_2692[0:0];
  _RAND_2693 = {1{`RANDOM}};
  mesh_0_12_io_in_control_1_propagate_pipe_b = _RAND_2693[0:0];
  _RAND_2694 = {1{`RANDOM}};
  mesh_1_12_io_in_control_0_shift_pipe_b = _RAND_2694[4:0];
  _RAND_2695 = {1{`RANDOM}};
  mesh_1_12_io_in_control_0_dataflow_pipe_b = _RAND_2695[0:0];
  _RAND_2696 = {1{`RANDOM}};
  mesh_1_12_io_in_control_0_propagate_pipe_b = _RAND_2696[0:0];
  _RAND_2697 = {1{`RANDOM}};
  mesh_1_12_io_in_control_1_shift_pipe_b = _RAND_2697[4:0];
  _RAND_2698 = {1{`RANDOM}};
  mesh_1_12_io_in_control_1_dataflow_pipe_b = _RAND_2698[0:0];
  _RAND_2699 = {1{`RANDOM}};
  mesh_1_12_io_in_control_1_propagate_pipe_b = _RAND_2699[0:0];
  _RAND_2700 = {1{`RANDOM}};
  mesh_2_12_io_in_control_0_shift_pipe_b = _RAND_2700[4:0];
  _RAND_2701 = {1{`RANDOM}};
  mesh_2_12_io_in_control_0_dataflow_pipe_b = _RAND_2701[0:0];
  _RAND_2702 = {1{`RANDOM}};
  mesh_2_12_io_in_control_0_propagate_pipe_b = _RAND_2702[0:0];
  _RAND_2703 = {1{`RANDOM}};
  mesh_2_12_io_in_control_1_shift_pipe_b = _RAND_2703[4:0];
  _RAND_2704 = {1{`RANDOM}};
  mesh_2_12_io_in_control_1_dataflow_pipe_b = _RAND_2704[0:0];
  _RAND_2705 = {1{`RANDOM}};
  mesh_2_12_io_in_control_1_propagate_pipe_b = _RAND_2705[0:0];
  _RAND_2706 = {1{`RANDOM}};
  mesh_3_12_io_in_control_0_shift_pipe_b = _RAND_2706[4:0];
  _RAND_2707 = {1{`RANDOM}};
  mesh_3_12_io_in_control_0_dataflow_pipe_b = _RAND_2707[0:0];
  _RAND_2708 = {1{`RANDOM}};
  mesh_3_12_io_in_control_0_propagate_pipe_b = _RAND_2708[0:0];
  _RAND_2709 = {1{`RANDOM}};
  mesh_3_12_io_in_control_1_shift_pipe_b = _RAND_2709[4:0];
  _RAND_2710 = {1{`RANDOM}};
  mesh_3_12_io_in_control_1_dataflow_pipe_b = _RAND_2710[0:0];
  _RAND_2711 = {1{`RANDOM}};
  mesh_3_12_io_in_control_1_propagate_pipe_b = _RAND_2711[0:0];
  _RAND_2712 = {1{`RANDOM}};
  mesh_4_12_io_in_control_0_shift_pipe_b = _RAND_2712[4:0];
  _RAND_2713 = {1{`RANDOM}};
  mesh_4_12_io_in_control_0_dataflow_pipe_b = _RAND_2713[0:0];
  _RAND_2714 = {1{`RANDOM}};
  mesh_4_12_io_in_control_0_propagate_pipe_b = _RAND_2714[0:0];
  _RAND_2715 = {1{`RANDOM}};
  mesh_4_12_io_in_control_1_shift_pipe_b = _RAND_2715[4:0];
  _RAND_2716 = {1{`RANDOM}};
  mesh_4_12_io_in_control_1_dataflow_pipe_b = _RAND_2716[0:0];
  _RAND_2717 = {1{`RANDOM}};
  mesh_4_12_io_in_control_1_propagate_pipe_b = _RAND_2717[0:0];
  _RAND_2718 = {1{`RANDOM}};
  mesh_5_12_io_in_control_0_shift_pipe_b = _RAND_2718[4:0];
  _RAND_2719 = {1{`RANDOM}};
  mesh_5_12_io_in_control_0_dataflow_pipe_b = _RAND_2719[0:0];
  _RAND_2720 = {1{`RANDOM}};
  mesh_5_12_io_in_control_0_propagate_pipe_b = _RAND_2720[0:0];
  _RAND_2721 = {1{`RANDOM}};
  mesh_5_12_io_in_control_1_shift_pipe_b = _RAND_2721[4:0];
  _RAND_2722 = {1{`RANDOM}};
  mesh_5_12_io_in_control_1_dataflow_pipe_b = _RAND_2722[0:0];
  _RAND_2723 = {1{`RANDOM}};
  mesh_5_12_io_in_control_1_propagate_pipe_b = _RAND_2723[0:0];
  _RAND_2724 = {1{`RANDOM}};
  mesh_6_12_io_in_control_0_shift_pipe_b = _RAND_2724[4:0];
  _RAND_2725 = {1{`RANDOM}};
  mesh_6_12_io_in_control_0_dataflow_pipe_b = _RAND_2725[0:0];
  _RAND_2726 = {1{`RANDOM}};
  mesh_6_12_io_in_control_0_propagate_pipe_b = _RAND_2726[0:0];
  _RAND_2727 = {1{`RANDOM}};
  mesh_6_12_io_in_control_1_shift_pipe_b = _RAND_2727[4:0];
  _RAND_2728 = {1{`RANDOM}};
  mesh_6_12_io_in_control_1_dataflow_pipe_b = _RAND_2728[0:0];
  _RAND_2729 = {1{`RANDOM}};
  mesh_6_12_io_in_control_1_propagate_pipe_b = _RAND_2729[0:0];
  _RAND_2730 = {1{`RANDOM}};
  mesh_7_12_io_in_control_0_shift_pipe_b = _RAND_2730[4:0];
  _RAND_2731 = {1{`RANDOM}};
  mesh_7_12_io_in_control_0_dataflow_pipe_b = _RAND_2731[0:0];
  _RAND_2732 = {1{`RANDOM}};
  mesh_7_12_io_in_control_0_propagate_pipe_b = _RAND_2732[0:0];
  _RAND_2733 = {1{`RANDOM}};
  mesh_7_12_io_in_control_1_shift_pipe_b = _RAND_2733[4:0];
  _RAND_2734 = {1{`RANDOM}};
  mesh_7_12_io_in_control_1_dataflow_pipe_b = _RAND_2734[0:0];
  _RAND_2735 = {1{`RANDOM}};
  mesh_7_12_io_in_control_1_propagate_pipe_b = _RAND_2735[0:0];
  _RAND_2736 = {1{`RANDOM}};
  mesh_8_12_io_in_control_0_shift_pipe_b = _RAND_2736[4:0];
  _RAND_2737 = {1{`RANDOM}};
  mesh_8_12_io_in_control_0_dataflow_pipe_b = _RAND_2737[0:0];
  _RAND_2738 = {1{`RANDOM}};
  mesh_8_12_io_in_control_0_propagate_pipe_b = _RAND_2738[0:0];
  _RAND_2739 = {1{`RANDOM}};
  mesh_8_12_io_in_control_1_shift_pipe_b = _RAND_2739[4:0];
  _RAND_2740 = {1{`RANDOM}};
  mesh_8_12_io_in_control_1_dataflow_pipe_b = _RAND_2740[0:0];
  _RAND_2741 = {1{`RANDOM}};
  mesh_8_12_io_in_control_1_propagate_pipe_b = _RAND_2741[0:0];
  _RAND_2742 = {1{`RANDOM}};
  mesh_9_12_io_in_control_0_shift_pipe_b = _RAND_2742[4:0];
  _RAND_2743 = {1{`RANDOM}};
  mesh_9_12_io_in_control_0_dataflow_pipe_b = _RAND_2743[0:0];
  _RAND_2744 = {1{`RANDOM}};
  mesh_9_12_io_in_control_0_propagate_pipe_b = _RAND_2744[0:0];
  _RAND_2745 = {1{`RANDOM}};
  mesh_9_12_io_in_control_1_shift_pipe_b = _RAND_2745[4:0];
  _RAND_2746 = {1{`RANDOM}};
  mesh_9_12_io_in_control_1_dataflow_pipe_b = _RAND_2746[0:0];
  _RAND_2747 = {1{`RANDOM}};
  mesh_9_12_io_in_control_1_propagate_pipe_b = _RAND_2747[0:0];
  _RAND_2748 = {1{`RANDOM}};
  mesh_10_12_io_in_control_0_shift_pipe_b = _RAND_2748[4:0];
  _RAND_2749 = {1{`RANDOM}};
  mesh_10_12_io_in_control_0_dataflow_pipe_b = _RAND_2749[0:0];
  _RAND_2750 = {1{`RANDOM}};
  mesh_10_12_io_in_control_0_propagate_pipe_b = _RAND_2750[0:0];
  _RAND_2751 = {1{`RANDOM}};
  mesh_10_12_io_in_control_1_shift_pipe_b = _RAND_2751[4:0];
  _RAND_2752 = {1{`RANDOM}};
  mesh_10_12_io_in_control_1_dataflow_pipe_b = _RAND_2752[0:0];
  _RAND_2753 = {1{`RANDOM}};
  mesh_10_12_io_in_control_1_propagate_pipe_b = _RAND_2753[0:0];
  _RAND_2754 = {1{`RANDOM}};
  mesh_11_12_io_in_control_0_shift_pipe_b = _RAND_2754[4:0];
  _RAND_2755 = {1{`RANDOM}};
  mesh_11_12_io_in_control_0_dataflow_pipe_b = _RAND_2755[0:0];
  _RAND_2756 = {1{`RANDOM}};
  mesh_11_12_io_in_control_0_propagate_pipe_b = _RAND_2756[0:0];
  _RAND_2757 = {1{`RANDOM}};
  mesh_11_12_io_in_control_1_shift_pipe_b = _RAND_2757[4:0];
  _RAND_2758 = {1{`RANDOM}};
  mesh_11_12_io_in_control_1_dataflow_pipe_b = _RAND_2758[0:0];
  _RAND_2759 = {1{`RANDOM}};
  mesh_11_12_io_in_control_1_propagate_pipe_b = _RAND_2759[0:0];
  _RAND_2760 = {1{`RANDOM}};
  mesh_12_12_io_in_control_0_shift_pipe_b = _RAND_2760[4:0];
  _RAND_2761 = {1{`RANDOM}};
  mesh_12_12_io_in_control_0_dataflow_pipe_b = _RAND_2761[0:0];
  _RAND_2762 = {1{`RANDOM}};
  mesh_12_12_io_in_control_0_propagate_pipe_b = _RAND_2762[0:0];
  _RAND_2763 = {1{`RANDOM}};
  mesh_12_12_io_in_control_1_shift_pipe_b = _RAND_2763[4:0];
  _RAND_2764 = {1{`RANDOM}};
  mesh_12_12_io_in_control_1_dataflow_pipe_b = _RAND_2764[0:0];
  _RAND_2765 = {1{`RANDOM}};
  mesh_12_12_io_in_control_1_propagate_pipe_b = _RAND_2765[0:0];
  _RAND_2766 = {1{`RANDOM}};
  mesh_13_12_io_in_control_0_shift_pipe_b = _RAND_2766[4:0];
  _RAND_2767 = {1{`RANDOM}};
  mesh_13_12_io_in_control_0_dataflow_pipe_b = _RAND_2767[0:0];
  _RAND_2768 = {1{`RANDOM}};
  mesh_13_12_io_in_control_0_propagate_pipe_b = _RAND_2768[0:0];
  _RAND_2769 = {1{`RANDOM}};
  mesh_13_12_io_in_control_1_shift_pipe_b = _RAND_2769[4:0];
  _RAND_2770 = {1{`RANDOM}};
  mesh_13_12_io_in_control_1_dataflow_pipe_b = _RAND_2770[0:0];
  _RAND_2771 = {1{`RANDOM}};
  mesh_13_12_io_in_control_1_propagate_pipe_b = _RAND_2771[0:0];
  _RAND_2772 = {1{`RANDOM}};
  mesh_14_12_io_in_control_0_shift_pipe_b = _RAND_2772[4:0];
  _RAND_2773 = {1{`RANDOM}};
  mesh_14_12_io_in_control_0_dataflow_pipe_b = _RAND_2773[0:0];
  _RAND_2774 = {1{`RANDOM}};
  mesh_14_12_io_in_control_0_propagate_pipe_b = _RAND_2774[0:0];
  _RAND_2775 = {1{`RANDOM}};
  mesh_14_12_io_in_control_1_shift_pipe_b = _RAND_2775[4:0];
  _RAND_2776 = {1{`RANDOM}};
  mesh_14_12_io_in_control_1_dataflow_pipe_b = _RAND_2776[0:0];
  _RAND_2777 = {1{`RANDOM}};
  mesh_14_12_io_in_control_1_propagate_pipe_b = _RAND_2777[0:0];
  _RAND_2778 = {1{`RANDOM}};
  mesh_15_12_io_in_control_0_shift_pipe_b = _RAND_2778[4:0];
  _RAND_2779 = {1{`RANDOM}};
  mesh_15_12_io_in_control_0_dataflow_pipe_b = _RAND_2779[0:0];
  _RAND_2780 = {1{`RANDOM}};
  mesh_15_12_io_in_control_0_propagate_pipe_b = _RAND_2780[0:0];
  _RAND_2781 = {1{`RANDOM}};
  mesh_15_12_io_in_control_1_shift_pipe_b = _RAND_2781[4:0];
  _RAND_2782 = {1{`RANDOM}};
  mesh_15_12_io_in_control_1_dataflow_pipe_b = _RAND_2782[0:0];
  _RAND_2783 = {1{`RANDOM}};
  mesh_15_12_io_in_control_1_propagate_pipe_b = _RAND_2783[0:0];
  _RAND_2784 = {1{`RANDOM}};
  mesh_0_13_io_in_control_0_shift_pipe_b = _RAND_2784[4:0];
  _RAND_2785 = {1{`RANDOM}};
  mesh_0_13_io_in_control_0_dataflow_pipe_b = _RAND_2785[0:0];
  _RAND_2786 = {1{`RANDOM}};
  mesh_0_13_io_in_control_0_propagate_pipe_b = _RAND_2786[0:0];
  _RAND_2787 = {1{`RANDOM}};
  mesh_0_13_io_in_control_1_shift_pipe_b = _RAND_2787[4:0];
  _RAND_2788 = {1{`RANDOM}};
  mesh_0_13_io_in_control_1_dataflow_pipe_b = _RAND_2788[0:0];
  _RAND_2789 = {1{`RANDOM}};
  mesh_0_13_io_in_control_1_propagate_pipe_b = _RAND_2789[0:0];
  _RAND_2790 = {1{`RANDOM}};
  mesh_1_13_io_in_control_0_shift_pipe_b = _RAND_2790[4:0];
  _RAND_2791 = {1{`RANDOM}};
  mesh_1_13_io_in_control_0_dataflow_pipe_b = _RAND_2791[0:0];
  _RAND_2792 = {1{`RANDOM}};
  mesh_1_13_io_in_control_0_propagate_pipe_b = _RAND_2792[0:0];
  _RAND_2793 = {1{`RANDOM}};
  mesh_1_13_io_in_control_1_shift_pipe_b = _RAND_2793[4:0];
  _RAND_2794 = {1{`RANDOM}};
  mesh_1_13_io_in_control_1_dataflow_pipe_b = _RAND_2794[0:0];
  _RAND_2795 = {1{`RANDOM}};
  mesh_1_13_io_in_control_1_propagate_pipe_b = _RAND_2795[0:0];
  _RAND_2796 = {1{`RANDOM}};
  mesh_2_13_io_in_control_0_shift_pipe_b = _RAND_2796[4:0];
  _RAND_2797 = {1{`RANDOM}};
  mesh_2_13_io_in_control_0_dataflow_pipe_b = _RAND_2797[0:0];
  _RAND_2798 = {1{`RANDOM}};
  mesh_2_13_io_in_control_0_propagate_pipe_b = _RAND_2798[0:0];
  _RAND_2799 = {1{`RANDOM}};
  mesh_2_13_io_in_control_1_shift_pipe_b = _RAND_2799[4:0];
  _RAND_2800 = {1{`RANDOM}};
  mesh_2_13_io_in_control_1_dataflow_pipe_b = _RAND_2800[0:0];
  _RAND_2801 = {1{`RANDOM}};
  mesh_2_13_io_in_control_1_propagate_pipe_b = _RAND_2801[0:0];
  _RAND_2802 = {1{`RANDOM}};
  mesh_3_13_io_in_control_0_shift_pipe_b = _RAND_2802[4:0];
  _RAND_2803 = {1{`RANDOM}};
  mesh_3_13_io_in_control_0_dataflow_pipe_b = _RAND_2803[0:0];
  _RAND_2804 = {1{`RANDOM}};
  mesh_3_13_io_in_control_0_propagate_pipe_b = _RAND_2804[0:0];
  _RAND_2805 = {1{`RANDOM}};
  mesh_3_13_io_in_control_1_shift_pipe_b = _RAND_2805[4:0];
  _RAND_2806 = {1{`RANDOM}};
  mesh_3_13_io_in_control_1_dataflow_pipe_b = _RAND_2806[0:0];
  _RAND_2807 = {1{`RANDOM}};
  mesh_3_13_io_in_control_1_propagate_pipe_b = _RAND_2807[0:0];
  _RAND_2808 = {1{`RANDOM}};
  mesh_4_13_io_in_control_0_shift_pipe_b = _RAND_2808[4:0];
  _RAND_2809 = {1{`RANDOM}};
  mesh_4_13_io_in_control_0_dataflow_pipe_b = _RAND_2809[0:0];
  _RAND_2810 = {1{`RANDOM}};
  mesh_4_13_io_in_control_0_propagate_pipe_b = _RAND_2810[0:0];
  _RAND_2811 = {1{`RANDOM}};
  mesh_4_13_io_in_control_1_shift_pipe_b = _RAND_2811[4:0];
  _RAND_2812 = {1{`RANDOM}};
  mesh_4_13_io_in_control_1_dataflow_pipe_b = _RAND_2812[0:0];
  _RAND_2813 = {1{`RANDOM}};
  mesh_4_13_io_in_control_1_propagate_pipe_b = _RAND_2813[0:0];
  _RAND_2814 = {1{`RANDOM}};
  mesh_5_13_io_in_control_0_shift_pipe_b = _RAND_2814[4:0];
  _RAND_2815 = {1{`RANDOM}};
  mesh_5_13_io_in_control_0_dataflow_pipe_b = _RAND_2815[0:0];
  _RAND_2816 = {1{`RANDOM}};
  mesh_5_13_io_in_control_0_propagate_pipe_b = _RAND_2816[0:0];
  _RAND_2817 = {1{`RANDOM}};
  mesh_5_13_io_in_control_1_shift_pipe_b = _RAND_2817[4:0];
  _RAND_2818 = {1{`RANDOM}};
  mesh_5_13_io_in_control_1_dataflow_pipe_b = _RAND_2818[0:0];
  _RAND_2819 = {1{`RANDOM}};
  mesh_5_13_io_in_control_1_propagate_pipe_b = _RAND_2819[0:0];
  _RAND_2820 = {1{`RANDOM}};
  mesh_6_13_io_in_control_0_shift_pipe_b = _RAND_2820[4:0];
  _RAND_2821 = {1{`RANDOM}};
  mesh_6_13_io_in_control_0_dataflow_pipe_b = _RAND_2821[0:0];
  _RAND_2822 = {1{`RANDOM}};
  mesh_6_13_io_in_control_0_propagate_pipe_b = _RAND_2822[0:0];
  _RAND_2823 = {1{`RANDOM}};
  mesh_6_13_io_in_control_1_shift_pipe_b = _RAND_2823[4:0];
  _RAND_2824 = {1{`RANDOM}};
  mesh_6_13_io_in_control_1_dataflow_pipe_b = _RAND_2824[0:0];
  _RAND_2825 = {1{`RANDOM}};
  mesh_6_13_io_in_control_1_propagate_pipe_b = _RAND_2825[0:0];
  _RAND_2826 = {1{`RANDOM}};
  mesh_7_13_io_in_control_0_shift_pipe_b = _RAND_2826[4:0];
  _RAND_2827 = {1{`RANDOM}};
  mesh_7_13_io_in_control_0_dataflow_pipe_b = _RAND_2827[0:0];
  _RAND_2828 = {1{`RANDOM}};
  mesh_7_13_io_in_control_0_propagate_pipe_b = _RAND_2828[0:0];
  _RAND_2829 = {1{`RANDOM}};
  mesh_7_13_io_in_control_1_shift_pipe_b = _RAND_2829[4:0];
  _RAND_2830 = {1{`RANDOM}};
  mesh_7_13_io_in_control_1_dataflow_pipe_b = _RAND_2830[0:0];
  _RAND_2831 = {1{`RANDOM}};
  mesh_7_13_io_in_control_1_propagate_pipe_b = _RAND_2831[0:0];
  _RAND_2832 = {1{`RANDOM}};
  mesh_8_13_io_in_control_0_shift_pipe_b = _RAND_2832[4:0];
  _RAND_2833 = {1{`RANDOM}};
  mesh_8_13_io_in_control_0_dataflow_pipe_b = _RAND_2833[0:0];
  _RAND_2834 = {1{`RANDOM}};
  mesh_8_13_io_in_control_0_propagate_pipe_b = _RAND_2834[0:0];
  _RAND_2835 = {1{`RANDOM}};
  mesh_8_13_io_in_control_1_shift_pipe_b = _RAND_2835[4:0];
  _RAND_2836 = {1{`RANDOM}};
  mesh_8_13_io_in_control_1_dataflow_pipe_b = _RAND_2836[0:0];
  _RAND_2837 = {1{`RANDOM}};
  mesh_8_13_io_in_control_1_propagate_pipe_b = _RAND_2837[0:0];
  _RAND_2838 = {1{`RANDOM}};
  mesh_9_13_io_in_control_0_shift_pipe_b = _RAND_2838[4:0];
  _RAND_2839 = {1{`RANDOM}};
  mesh_9_13_io_in_control_0_dataflow_pipe_b = _RAND_2839[0:0];
  _RAND_2840 = {1{`RANDOM}};
  mesh_9_13_io_in_control_0_propagate_pipe_b = _RAND_2840[0:0];
  _RAND_2841 = {1{`RANDOM}};
  mesh_9_13_io_in_control_1_shift_pipe_b = _RAND_2841[4:0];
  _RAND_2842 = {1{`RANDOM}};
  mesh_9_13_io_in_control_1_dataflow_pipe_b = _RAND_2842[0:0];
  _RAND_2843 = {1{`RANDOM}};
  mesh_9_13_io_in_control_1_propagate_pipe_b = _RAND_2843[0:0];
  _RAND_2844 = {1{`RANDOM}};
  mesh_10_13_io_in_control_0_shift_pipe_b = _RAND_2844[4:0];
  _RAND_2845 = {1{`RANDOM}};
  mesh_10_13_io_in_control_0_dataflow_pipe_b = _RAND_2845[0:0];
  _RAND_2846 = {1{`RANDOM}};
  mesh_10_13_io_in_control_0_propagate_pipe_b = _RAND_2846[0:0];
  _RAND_2847 = {1{`RANDOM}};
  mesh_10_13_io_in_control_1_shift_pipe_b = _RAND_2847[4:0];
  _RAND_2848 = {1{`RANDOM}};
  mesh_10_13_io_in_control_1_dataflow_pipe_b = _RAND_2848[0:0];
  _RAND_2849 = {1{`RANDOM}};
  mesh_10_13_io_in_control_1_propagate_pipe_b = _RAND_2849[0:0];
  _RAND_2850 = {1{`RANDOM}};
  mesh_11_13_io_in_control_0_shift_pipe_b = _RAND_2850[4:0];
  _RAND_2851 = {1{`RANDOM}};
  mesh_11_13_io_in_control_0_dataflow_pipe_b = _RAND_2851[0:0];
  _RAND_2852 = {1{`RANDOM}};
  mesh_11_13_io_in_control_0_propagate_pipe_b = _RAND_2852[0:0];
  _RAND_2853 = {1{`RANDOM}};
  mesh_11_13_io_in_control_1_shift_pipe_b = _RAND_2853[4:0];
  _RAND_2854 = {1{`RANDOM}};
  mesh_11_13_io_in_control_1_dataflow_pipe_b = _RAND_2854[0:0];
  _RAND_2855 = {1{`RANDOM}};
  mesh_11_13_io_in_control_1_propagate_pipe_b = _RAND_2855[0:0];
  _RAND_2856 = {1{`RANDOM}};
  mesh_12_13_io_in_control_0_shift_pipe_b = _RAND_2856[4:0];
  _RAND_2857 = {1{`RANDOM}};
  mesh_12_13_io_in_control_0_dataflow_pipe_b = _RAND_2857[0:0];
  _RAND_2858 = {1{`RANDOM}};
  mesh_12_13_io_in_control_0_propagate_pipe_b = _RAND_2858[0:0];
  _RAND_2859 = {1{`RANDOM}};
  mesh_12_13_io_in_control_1_shift_pipe_b = _RAND_2859[4:0];
  _RAND_2860 = {1{`RANDOM}};
  mesh_12_13_io_in_control_1_dataflow_pipe_b = _RAND_2860[0:0];
  _RAND_2861 = {1{`RANDOM}};
  mesh_12_13_io_in_control_1_propagate_pipe_b = _RAND_2861[0:0];
  _RAND_2862 = {1{`RANDOM}};
  mesh_13_13_io_in_control_0_shift_pipe_b = _RAND_2862[4:0];
  _RAND_2863 = {1{`RANDOM}};
  mesh_13_13_io_in_control_0_dataflow_pipe_b = _RAND_2863[0:0];
  _RAND_2864 = {1{`RANDOM}};
  mesh_13_13_io_in_control_0_propagate_pipe_b = _RAND_2864[0:0];
  _RAND_2865 = {1{`RANDOM}};
  mesh_13_13_io_in_control_1_shift_pipe_b = _RAND_2865[4:0];
  _RAND_2866 = {1{`RANDOM}};
  mesh_13_13_io_in_control_1_dataflow_pipe_b = _RAND_2866[0:0];
  _RAND_2867 = {1{`RANDOM}};
  mesh_13_13_io_in_control_1_propagate_pipe_b = _RAND_2867[0:0];
  _RAND_2868 = {1{`RANDOM}};
  mesh_14_13_io_in_control_0_shift_pipe_b = _RAND_2868[4:0];
  _RAND_2869 = {1{`RANDOM}};
  mesh_14_13_io_in_control_0_dataflow_pipe_b = _RAND_2869[0:0];
  _RAND_2870 = {1{`RANDOM}};
  mesh_14_13_io_in_control_0_propagate_pipe_b = _RAND_2870[0:0];
  _RAND_2871 = {1{`RANDOM}};
  mesh_14_13_io_in_control_1_shift_pipe_b = _RAND_2871[4:0];
  _RAND_2872 = {1{`RANDOM}};
  mesh_14_13_io_in_control_1_dataflow_pipe_b = _RAND_2872[0:0];
  _RAND_2873 = {1{`RANDOM}};
  mesh_14_13_io_in_control_1_propagate_pipe_b = _RAND_2873[0:0];
  _RAND_2874 = {1{`RANDOM}};
  mesh_15_13_io_in_control_0_shift_pipe_b = _RAND_2874[4:0];
  _RAND_2875 = {1{`RANDOM}};
  mesh_15_13_io_in_control_0_dataflow_pipe_b = _RAND_2875[0:0];
  _RAND_2876 = {1{`RANDOM}};
  mesh_15_13_io_in_control_0_propagate_pipe_b = _RAND_2876[0:0];
  _RAND_2877 = {1{`RANDOM}};
  mesh_15_13_io_in_control_1_shift_pipe_b = _RAND_2877[4:0];
  _RAND_2878 = {1{`RANDOM}};
  mesh_15_13_io_in_control_1_dataflow_pipe_b = _RAND_2878[0:0];
  _RAND_2879 = {1{`RANDOM}};
  mesh_15_13_io_in_control_1_propagate_pipe_b = _RAND_2879[0:0];
  _RAND_2880 = {1{`RANDOM}};
  mesh_0_14_io_in_control_0_shift_pipe_b = _RAND_2880[4:0];
  _RAND_2881 = {1{`RANDOM}};
  mesh_0_14_io_in_control_0_dataflow_pipe_b = _RAND_2881[0:0];
  _RAND_2882 = {1{`RANDOM}};
  mesh_0_14_io_in_control_0_propagate_pipe_b = _RAND_2882[0:0];
  _RAND_2883 = {1{`RANDOM}};
  mesh_0_14_io_in_control_1_shift_pipe_b = _RAND_2883[4:0];
  _RAND_2884 = {1{`RANDOM}};
  mesh_0_14_io_in_control_1_dataflow_pipe_b = _RAND_2884[0:0];
  _RAND_2885 = {1{`RANDOM}};
  mesh_0_14_io_in_control_1_propagate_pipe_b = _RAND_2885[0:0];
  _RAND_2886 = {1{`RANDOM}};
  mesh_1_14_io_in_control_0_shift_pipe_b = _RAND_2886[4:0];
  _RAND_2887 = {1{`RANDOM}};
  mesh_1_14_io_in_control_0_dataflow_pipe_b = _RAND_2887[0:0];
  _RAND_2888 = {1{`RANDOM}};
  mesh_1_14_io_in_control_0_propagate_pipe_b = _RAND_2888[0:0];
  _RAND_2889 = {1{`RANDOM}};
  mesh_1_14_io_in_control_1_shift_pipe_b = _RAND_2889[4:0];
  _RAND_2890 = {1{`RANDOM}};
  mesh_1_14_io_in_control_1_dataflow_pipe_b = _RAND_2890[0:0];
  _RAND_2891 = {1{`RANDOM}};
  mesh_1_14_io_in_control_1_propagate_pipe_b = _RAND_2891[0:0];
  _RAND_2892 = {1{`RANDOM}};
  mesh_2_14_io_in_control_0_shift_pipe_b = _RAND_2892[4:0];
  _RAND_2893 = {1{`RANDOM}};
  mesh_2_14_io_in_control_0_dataflow_pipe_b = _RAND_2893[0:0];
  _RAND_2894 = {1{`RANDOM}};
  mesh_2_14_io_in_control_0_propagate_pipe_b = _RAND_2894[0:0];
  _RAND_2895 = {1{`RANDOM}};
  mesh_2_14_io_in_control_1_shift_pipe_b = _RAND_2895[4:0];
  _RAND_2896 = {1{`RANDOM}};
  mesh_2_14_io_in_control_1_dataflow_pipe_b = _RAND_2896[0:0];
  _RAND_2897 = {1{`RANDOM}};
  mesh_2_14_io_in_control_1_propagate_pipe_b = _RAND_2897[0:0];
  _RAND_2898 = {1{`RANDOM}};
  mesh_3_14_io_in_control_0_shift_pipe_b = _RAND_2898[4:0];
  _RAND_2899 = {1{`RANDOM}};
  mesh_3_14_io_in_control_0_dataflow_pipe_b = _RAND_2899[0:0];
  _RAND_2900 = {1{`RANDOM}};
  mesh_3_14_io_in_control_0_propagate_pipe_b = _RAND_2900[0:0];
  _RAND_2901 = {1{`RANDOM}};
  mesh_3_14_io_in_control_1_shift_pipe_b = _RAND_2901[4:0];
  _RAND_2902 = {1{`RANDOM}};
  mesh_3_14_io_in_control_1_dataflow_pipe_b = _RAND_2902[0:0];
  _RAND_2903 = {1{`RANDOM}};
  mesh_3_14_io_in_control_1_propagate_pipe_b = _RAND_2903[0:0];
  _RAND_2904 = {1{`RANDOM}};
  mesh_4_14_io_in_control_0_shift_pipe_b = _RAND_2904[4:0];
  _RAND_2905 = {1{`RANDOM}};
  mesh_4_14_io_in_control_0_dataflow_pipe_b = _RAND_2905[0:0];
  _RAND_2906 = {1{`RANDOM}};
  mesh_4_14_io_in_control_0_propagate_pipe_b = _RAND_2906[0:0];
  _RAND_2907 = {1{`RANDOM}};
  mesh_4_14_io_in_control_1_shift_pipe_b = _RAND_2907[4:0];
  _RAND_2908 = {1{`RANDOM}};
  mesh_4_14_io_in_control_1_dataflow_pipe_b = _RAND_2908[0:0];
  _RAND_2909 = {1{`RANDOM}};
  mesh_4_14_io_in_control_1_propagate_pipe_b = _RAND_2909[0:0];
  _RAND_2910 = {1{`RANDOM}};
  mesh_5_14_io_in_control_0_shift_pipe_b = _RAND_2910[4:0];
  _RAND_2911 = {1{`RANDOM}};
  mesh_5_14_io_in_control_0_dataflow_pipe_b = _RAND_2911[0:0];
  _RAND_2912 = {1{`RANDOM}};
  mesh_5_14_io_in_control_0_propagate_pipe_b = _RAND_2912[0:0];
  _RAND_2913 = {1{`RANDOM}};
  mesh_5_14_io_in_control_1_shift_pipe_b = _RAND_2913[4:0];
  _RAND_2914 = {1{`RANDOM}};
  mesh_5_14_io_in_control_1_dataflow_pipe_b = _RAND_2914[0:0];
  _RAND_2915 = {1{`RANDOM}};
  mesh_5_14_io_in_control_1_propagate_pipe_b = _RAND_2915[0:0];
  _RAND_2916 = {1{`RANDOM}};
  mesh_6_14_io_in_control_0_shift_pipe_b = _RAND_2916[4:0];
  _RAND_2917 = {1{`RANDOM}};
  mesh_6_14_io_in_control_0_dataflow_pipe_b = _RAND_2917[0:0];
  _RAND_2918 = {1{`RANDOM}};
  mesh_6_14_io_in_control_0_propagate_pipe_b = _RAND_2918[0:0];
  _RAND_2919 = {1{`RANDOM}};
  mesh_6_14_io_in_control_1_shift_pipe_b = _RAND_2919[4:0];
  _RAND_2920 = {1{`RANDOM}};
  mesh_6_14_io_in_control_1_dataflow_pipe_b = _RAND_2920[0:0];
  _RAND_2921 = {1{`RANDOM}};
  mesh_6_14_io_in_control_1_propagate_pipe_b = _RAND_2921[0:0];
  _RAND_2922 = {1{`RANDOM}};
  mesh_7_14_io_in_control_0_shift_pipe_b = _RAND_2922[4:0];
  _RAND_2923 = {1{`RANDOM}};
  mesh_7_14_io_in_control_0_dataflow_pipe_b = _RAND_2923[0:0];
  _RAND_2924 = {1{`RANDOM}};
  mesh_7_14_io_in_control_0_propagate_pipe_b = _RAND_2924[0:0];
  _RAND_2925 = {1{`RANDOM}};
  mesh_7_14_io_in_control_1_shift_pipe_b = _RAND_2925[4:0];
  _RAND_2926 = {1{`RANDOM}};
  mesh_7_14_io_in_control_1_dataflow_pipe_b = _RAND_2926[0:0];
  _RAND_2927 = {1{`RANDOM}};
  mesh_7_14_io_in_control_1_propagate_pipe_b = _RAND_2927[0:0];
  _RAND_2928 = {1{`RANDOM}};
  mesh_8_14_io_in_control_0_shift_pipe_b = _RAND_2928[4:0];
  _RAND_2929 = {1{`RANDOM}};
  mesh_8_14_io_in_control_0_dataflow_pipe_b = _RAND_2929[0:0];
  _RAND_2930 = {1{`RANDOM}};
  mesh_8_14_io_in_control_0_propagate_pipe_b = _RAND_2930[0:0];
  _RAND_2931 = {1{`RANDOM}};
  mesh_8_14_io_in_control_1_shift_pipe_b = _RAND_2931[4:0];
  _RAND_2932 = {1{`RANDOM}};
  mesh_8_14_io_in_control_1_dataflow_pipe_b = _RAND_2932[0:0];
  _RAND_2933 = {1{`RANDOM}};
  mesh_8_14_io_in_control_1_propagate_pipe_b = _RAND_2933[0:0];
  _RAND_2934 = {1{`RANDOM}};
  mesh_9_14_io_in_control_0_shift_pipe_b = _RAND_2934[4:0];
  _RAND_2935 = {1{`RANDOM}};
  mesh_9_14_io_in_control_0_dataflow_pipe_b = _RAND_2935[0:0];
  _RAND_2936 = {1{`RANDOM}};
  mesh_9_14_io_in_control_0_propagate_pipe_b = _RAND_2936[0:0];
  _RAND_2937 = {1{`RANDOM}};
  mesh_9_14_io_in_control_1_shift_pipe_b = _RAND_2937[4:0];
  _RAND_2938 = {1{`RANDOM}};
  mesh_9_14_io_in_control_1_dataflow_pipe_b = _RAND_2938[0:0];
  _RAND_2939 = {1{`RANDOM}};
  mesh_9_14_io_in_control_1_propagate_pipe_b = _RAND_2939[0:0];
  _RAND_2940 = {1{`RANDOM}};
  mesh_10_14_io_in_control_0_shift_pipe_b = _RAND_2940[4:0];
  _RAND_2941 = {1{`RANDOM}};
  mesh_10_14_io_in_control_0_dataflow_pipe_b = _RAND_2941[0:0];
  _RAND_2942 = {1{`RANDOM}};
  mesh_10_14_io_in_control_0_propagate_pipe_b = _RAND_2942[0:0];
  _RAND_2943 = {1{`RANDOM}};
  mesh_10_14_io_in_control_1_shift_pipe_b = _RAND_2943[4:0];
  _RAND_2944 = {1{`RANDOM}};
  mesh_10_14_io_in_control_1_dataflow_pipe_b = _RAND_2944[0:0];
  _RAND_2945 = {1{`RANDOM}};
  mesh_10_14_io_in_control_1_propagate_pipe_b = _RAND_2945[0:0];
  _RAND_2946 = {1{`RANDOM}};
  mesh_11_14_io_in_control_0_shift_pipe_b = _RAND_2946[4:0];
  _RAND_2947 = {1{`RANDOM}};
  mesh_11_14_io_in_control_0_dataflow_pipe_b = _RAND_2947[0:0];
  _RAND_2948 = {1{`RANDOM}};
  mesh_11_14_io_in_control_0_propagate_pipe_b = _RAND_2948[0:0];
  _RAND_2949 = {1{`RANDOM}};
  mesh_11_14_io_in_control_1_shift_pipe_b = _RAND_2949[4:0];
  _RAND_2950 = {1{`RANDOM}};
  mesh_11_14_io_in_control_1_dataflow_pipe_b = _RAND_2950[0:0];
  _RAND_2951 = {1{`RANDOM}};
  mesh_11_14_io_in_control_1_propagate_pipe_b = _RAND_2951[0:0];
  _RAND_2952 = {1{`RANDOM}};
  mesh_12_14_io_in_control_0_shift_pipe_b = _RAND_2952[4:0];
  _RAND_2953 = {1{`RANDOM}};
  mesh_12_14_io_in_control_0_dataflow_pipe_b = _RAND_2953[0:0];
  _RAND_2954 = {1{`RANDOM}};
  mesh_12_14_io_in_control_0_propagate_pipe_b = _RAND_2954[0:0];
  _RAND_2955 = {1{`RANDOM}};
  mesh_12_14_io_in_control_1_shift_pipe_b = _RAND_2955[4:0];
  _RAND_2956 = {1{`RANDOM}};
  mesh_12_14_io_in_control_1_dataflow_pipe_b = _RAND_2956[0:0];
  _RAND_2957 = {1{`RANDOM}};
  mesh_12_14_io_in_control_1_propagate_pipe_b = _RAND_2957[0:0];
  _RAND_2958 = {1{`RANDOM}};
  mesh_13_14_io_in_control_0_shift_pipe_b = _RAND_2958[4:0];
  _RAND_2959 = {1{`RANDOM}};
  mesh_13_14_io_in_control_0_dataflow_pipe_b = _RAND_2959[0:0];
  _RAND_2960 = {1{`RANDOM}};
  mesh_13_14_io_in_control_0_propagate_pipe_b = _RAND_2960[0:0];
  _RAND_2961 = {1{`RANDOM}};
  mesh_13_14_io_in_control_1_shift_pipe_b = _RAND_2961[4:0];
  _RAND_2962 = {1{`RANDOM}};
  mesh_13_14_io_in_control_1_dataflow_pipe_b = _RAND_2962[0:0];
  _RAND_2963 = {1{`RANDOM}};
  mesh_13_14_io_in_control_1_propagate_pipe_b = _RAND_2963[0:0];
  _RAND_2964 = {1{`RANDOM}};
  mesh_14_14_io_in_control_0_shift_pipe_b = _RAND_2964[4:0];
  _RAND_2965 = {1{`RANDOM}};
  mesh_14_14_io_in_control_0_dataflow_pipe_b = _RAND_2965[0:0];
  _RAND_2966 = {1{`RANDOM}};
  mesh_14_14_io_in_control_0_propagate_pipe_b = _RAND_2966[0:0];
  _RAND_2967 = {1{`RANDOM}};
  mesh_14_14_io_in_control_1_shift_pipe_b = _RAND_2967[4:0];
  _RAND_2968 = {1{`RANDOM}};
  mesh_14_14_io_in_control_1_dataflow_pipe_b = _RAND_2968[0:0];
  _RAND_2969 = {1{`RANDOM}};
  mesh_14_14_io_in_control_1_propagate_pipe_b = _RAND_2969[0:0];
  _RAND_2970 = {1{`RANDOM}};
  mesh_15_14_io_in_control_0_shift_pipe_b = _RAND_2970[4:0];
  _RAND_2971 = {1{`RANDOM}};
  mesh_15_14_io_in_control_0_dataflow_pipe_b = _RAND_2971[0:0];
  _RAND_2972 = {1{`RANDOM}};
  mesh_15_14_io_in_control_0_propagate_pipe_b = _RAND_2972[0:0];
  _RAND_2973 = {1{`RANDOM}};
  mesh_15_14_io_in_control_1_shift_pipe_b = _RAND_2973[4:0];
  _RAND_2974 = {1{`RANDOM}};
  mesh_15_14_io_in_control_1_dataflow_pipe_b = _RAND_2974[0:0];
  _RAND_2975 = {1{`RANDOM}};
  mesh_15_14_io_in_control_1_propagate_pipe_b = _RAND_2975[0:0];
  _RAND_2976 = {1{`RANDOM}};
  mesh_0_15_io_in_control_0_shift_pipe_b = _RAND_2976[4:0];
  _RAND_2977 = {1{`RANDOM}};
  mesh_0_15_io_in_control_0_dataflow_pipe_b = _RAND_2977[0:0];
  _RAND_2978 = {1{`RANDOM}};
  mesh_0_15_io_in_control_0_propagate_pipe_b = _RAND_2978[0:0];
  _RAND_2979 = {1{`RANDOM}};
  mesh_0_15_io_in_control_1_shift_pipe_b = _RAND_2979[4:0];
  _RAND_2980 = {1{`RANDOM}};
  mesh_0_15_io_in_control_1_dataflow_pipe_b = _RAND_2980[0:0];
  _RAND_2981 = {1{`RANDOM}};
  mesh_0_15_io_in_control_1_propagate_pipe_b = _RAND_2981[0:0];
  _RAND_2982 = {1{`RANDOM}};
  mesh_1_15_io_in_control_0_shift_pipe_b = _RAND_2982[4:0];
  _RAND_2983 = {1{`RANDOM}};
  mesh_1_15_io_in_control_0_dataflow_pipe_b = _RAND_2983[0:0];
  _RAND_2984 = {1{`RANDOM}};
  mesh_1_15_io_in_control_0_propagate_pipe_b = _RAND_2984[0:0];
  _RAND_2985 = {1{`RANDOM}};
  mesh_1_15_io_in_control_1_shift_pipe_b = _RAND_2985[4:0];
  _RAND_2986 = {1{`RANDOM}};
  mesh_1_15_io_in_control_1_dataflow_pipe_b = _RAND_2986[0:0];
  _RAND_2987 = {1{`RANDOM}};
  mesh_1_15_io_in_control_1_propagate_pipe_b = _RAND_2987[0:0];
  _RAND_2988 = {1{`RANDOM}};
  mesh_2_15_io_in_control_0_shift_pipe_b = _RAND_2988[4:0];
  _RAND_2989 = {1{`RANDOM}};
  mesh_2_15_io_in_control_0_dataflow_pipe_b = _RAND_2989[0:0];
  _RAND_2990 = {1{`RANDOM}};
  mesh_2_15_io_in_control_0_propagate_pipe_b = _RAND_2990[0:0];
  _RAND_2991 = {1{`RANDOM}};
  mesh_2_15_io_in_control_1_shift_pipe_b = _RAND_2991[4:0];
  _RAND_2992 = {1{`RANDOM}};
  mesh_2_15_io_in_control_1_dataflow_pipe_b = _RAND_2992[0:0];
  _RAND_2993 = {1{`RANDOM}};
  mesh_2_15_io_in_control_1_propagate_pipe_b = _RAND_2993[0:0];
  _RAND_2994 = {1{`RANDOM}};
  mesh_3_15_io_in_control_0_shift_pipe_b = _RAND_2994[4:0];
  _RAND_2995 = {1{`RANDOM}};
  mesh_3_15_io_in_control_0_dataflow_pipe_b = _RAND_2995[0:0];
  _RAND_2996 = {1{`RANDOM}};
  mesh_3_15_io_in_control_0_propagate_pipe_b = _RAND_2996[0:0];
  _RAND_2997 = {1{`RANDOM}};
  mesh_3_15_io_in_control_1_shift_pipe_b = _RAND_2997[4:0];
  _RAND_2998 = {1{`RANDOM}};
  mesh_3_15_io_in_control_1_dataflow_pipe_b = _RAND_2998[0:0];
  _RAND_2999 = {1{`RANDOM}};
  mesh_3_15_io_in_control_1_propagate_pipe_b = _RAND_2999[0:0];
  _RAND_3000 = {1{`RANDOM}};
  mesh_4_15_io_in_control_0_shift_pipe_b = _RAND_3000[4:0];
  _RAND_3001 = {1{`RANDOM}};
  mesh_4_15_io_in_control_0_dataflow_pipe_b = _RAND_3001[0:0];
  _RAND_3002 = {1{`RANDOM}};
  mesh_4_15_io_in_control_0_propagate_pipe_b = _RAND_3002[0:0];
  _RAND_3003 = {1{`RANDOM}};
  mesh_4_15_io_in_control_1_shift_pipe_b = _RAND_3003[4:0];
  _RAND_3004 = {1{`RANDOM}};
  mesh_4_15_io_in_control_1_dataflow_pipe_b = _RAND_3004[0:0];
  _RAND_3005 = {1{`RANDOM}};
  mesh_4_15_io_in_control_1_propagate_pipe_b = _RAND_3005[0:0];
  _RAND_3006 = {1{`RANDOM}};
  mesh_5_15_io_in_control_0_shift_pipe_b = _RAND_3006[4:0];
  _RAND_3007 = {1{`RANDOM}};
  mesh_5_15_io_in_control_0_dataflow_pipe_b = _RAND_3007[0:0];
  _RAND_3008 = {1{`RANDOM}};
  mesh_5_15_io_in_control_0_propagate_pipe_b = _RAND_3008[0:0];
  _RAND_3009 = {1{`RANDOM}};
  mesh_5_15_io_in_control_1_shift_pipe_b = _RAND_3009[4:0];
  _RAND_3010 = {1{`RANDOM}};
  mesh_5_15_io_in_control_1_dataflow_pipe_b = _RAND_3010[0:0];
  _RAND_3011 = {1{`RANDOM}};
  mesh_5_15_io_in_control_1_propagate_pipe_b = _RAND_3011[0:0];
  _RAND_3012 = {1{`RANDOM}};
  mesh_6_15_io_in_control_0_shift_pipe_b = _RAND_3012[4:0];
  _RAND_3013 = {1{`RANDOM}};
  mesh_6_15_io_in_control_0_dataflow_pipe_b = _RAND_3013[0:0];
  _RAND_3014 = {1{`RANDOM}};
  mesh_6_15_io_in_control_0_propagate_pipe_b = _RAND_3014[0:0];
  _RAND_3015 = {1{`RANDOM}};
  mesh_6_15_io_in_control_1_shift_pipe_b = _RAND_3015[4:0];
  _RAND_3016 = {1{`RANDOM}};
  mesh_6_15_io_in_control_1_dataflow_pipe_b = _RAND_3016[0:0];
  _RAND_3017 = {1{`RANDOM}};
  mesh_6_15_io_in_control_1_propagate_pipe_b = _RAND_3017[0:0];
  _RAND_3018 = {1{`RANDOM}};
  mesh_7_15_io_in_control_0_shift_pipe_b = _RAND_3018[4:0];
  _RAND_3019 = {1{`RANDOM}};
  mesh_7_15_io_in_control_0_dataflow_pipe_b = _RAND_3019[0:0];
  _RAND_3020 = {1{`RANDOM}};
  mesh_7_15_io_in_control_0_propagate_pipe_b = _RAND_3020[0:0];
  _RAND_3021 = {1{`RANDOM}};
  mesh_7_15_io_in_control_1_shift_pipe_b = _RAND_3021[4:0];
  _RAND_3022 = {1{`RANDOM}};
  mesh_7_15_io_in_control_1_dataflow_pipe_b = _RAND_3022[0:0];
  _RAND_3023 = {1{`RANDOM}};
  mesh_7_15_io_in_control_1_propagate_pipe_b = _RAND_3023[0:0];
  _RAND_3024 = {1{`RANDOM}};
  mesh_8_15_io_in_control_0_shift_pipe_b = _RAND_3024[4:0];
  _RAND_3025 = {1{`RANDOM}};
  mesh_8_15_io_in_control_0_dataflow_pipe_b = _RAND_3025[0:0];
  _RAND_3026 = {1{`RANDOM}};
  mesh_8_15_io_in_control_0_propagate_pipe_b = _RAND_3026[0:0];
  _RAND_3027 = {1{`RANDOM}};
  mesh_8_15_io_in_control_1_shift_pipe_b = _RAND_3027[4:0];
  _RAND_3028 = {1{`RANDOM}};
  mesh_8_15_io_in_control_1_dataflow_pipe_b = _RAND_3028[0:0];
  _RAND_3029 = {1{`RANDOM}};
  mesh_8_15_io_in_control_1_propagate_pipe_b = _RAND_3029[0:0];
  _RAND_3030 = {1{`RANDOM}};
  mesh_9_15_io_in_control_0_shift_pipe_b = _RAND_3030[4:0];
  _RAND_3031 = {1{`RANDOM}};
  mesh_9_15_io_in_control_0_dataflow_pipe_b = _RAND_3031[0:0];
  _RAND_3032 = {1{`RANDOM}};
  mesh_9_15_io_in_control_0_propagate_pipe_b = _RAND_3032[0:0];
  _RAND_3033 = {1{`RANDOM}};
  mesh_9_15_io_in_control_1_shift_pipe_b = _RAND_3033[4:0];
  _RAND_3034 = {1{`RANDOM}};
  mesh_9_15_io_in_control_1_dataflow_pipe_b = _RAND_3034[0:0];
  _RAND_3035 = {1{`RANDOM}};
  mesh_9_15_io_in_control_1_propagate_pipe_b = _RAND_3035[0:0];
  _RAND_3036 = {1{`RANDOM}};
  mesh_10_15_io_in_control_0_shift_pipe_b = _RAND_3036[4:0];
  _RAND_3037 = {1{`RANDOM}};
  mesh_10_15_io_in_control_0_dataflow_pipe_b = _RAND_3037[0:0];
  _RAND_3038 = {1{`RANDOM}};
  mesh_10_15_io_in_control_0_propagate_pipe_b = _RAND_3038[0:0];
  _RAND_3039 = {1{`RANDOM}};
  mesh_10_15_io_in_control_1_shift_pipe_b = _RAND_3039[4:0];
  _RAND_3040 = {1{`RANDOM}};
  mesh_10_15_io_in_control_1_dataflow_pipe_b = _RAND_3040[0:0];
  _RAND_3041 = {1{`RANDOM}};
  mesh_10_15_io_in_control_1_propagate_pipe_b = _RAND_3041[0:0];
  _RAND_3042 = {1{`RANDOM}};
  mesh_11_15_io_in_control_0_shift_pipe_b = _RAND_3042[4:0];
  _RAND_3043 = {1{`RANDOM}};
  mesh_11_15_io_in_control_0_dataflow_pipe_b = _RAND_3043[0:0];
  _RAND_3044 = {1{`RANDOM}};
  mesh_11_15_io_in_control_0_propagate_pipe_b = _RAND_3044[0:0];
  _RAND_3045 = {1{`RANDOM}};
  mesh_11_15_io_in_control_1_shift_pipe_b = _RAND_3045[4:0];
  _RAND_3046 = {1{`RANDOM}};
  mesh_11_15_io_in_control_1_dataflow_pipe_b = _RAND_3046[0:0];
  _RAND_3047 = {1{`RANDOM}};
  mesh_11_15_io_in_control_1_propagate_pipe_b = _RAND_3047[0:0];
  _RAND_3048 = {1{`RANDOM}};
  mesh_12_15_io_in_control_0_shift_pipe_b = _RAND_3048[4:0];
  _RAND_3049 = {1{`RANDOM}};
  mesh_12_15_io_in_control_0_dataflow_pipe_b = _RAND_3049[0:0];
  _RAND_3050 = {1{`RANDOM}};
  mesh_12_15_io_in_control_0_propagate_pipe_b = _RAND_3050[0:0];
  _RAND_3051 = {1{`RANDOM}};
  mesh_12_15_io_in_control_1_shift_pipe_b = _RAND_3051[4:0];
  _RAND_3052 = {1{`RANDOM}};
  mesh_12_15_io_in_control_1_dataflow_pipe_b = _RAND_3052[0:0];
  _RAND_3053 = {1{`RANDOM}};
  mesh_12_15_io_in_control_1_propagate_pipe_b = _RAND_3053[0:0];
  _RAND_3054 = {1{`RANDOM}};
  mesh_13_15_io_in_control_0_shift_pipe_b = _RAND_3054[4:0];
  _RAND_3055 = {1{`RANDOM}};
  mesh_13_15_io_in_control_0_dataflow_pipe_b = _RAND_3055[0:0];
  _RAND_3056 = {1{`RANDOM}};
  mesh_13_15_io_in_control_0_propagate_pipe_b = _RAND_3056[0:0];
  _RAND_3057 = {1{`RANDOM}};
  mesh_13_15_io_in_control_1_shift_pipe_b = _RAND_3057[4:0];
  _RAND_3058 = {1{`RANDOM}};
  mesh_13_15_io_in_control_1_dataflow_pipe_b = _RAND_3058[0:0];
  _RAND_3059 = {1{`RANDOM}};
  mesh_13_15_io_in_control_1_propagate_pipe_b = _RAND_3059[0:0];
  _RAND_3060 = {1{`RANDOM}};
  mesh_14_15_io_in_control_0_shift_pipe_b = _RAND_3060[4:0];
  _RAND_3061 = {1{`RANDOM}};
  mesh_14_15_io_in_control_0_dataflow_pipe_b = _RAND_3061[0:0];
  _RAND_3062 = {1{`RANDOM}};
  mesh_14_15_io_in_control_0_propagate_pipe_b = _RAND_3062[0:0];
  _RAND_3063 = {1{`RANDOM}};
  mesh_14_15_io_in_control_1_shift_pipe_b = _RAND_3063[4:0];
  _RAND_3064 = {1{`RANDOM}};
  mesh_14_15_io_in_control_1_dataflow_pipe_b = _RAND_3064[0:0];
  _RAND_3065 = {1{`RANDOM}};
  mesh_14_15_io_in_control_1_propagate_pipe_b = _RAND_3065[0:0];
  _RAND_3066 = {1{`RANDOM}};
  mesh_15_15_io_in_control_0_shift_pipe_b = _RAND_3066[4:0];
  _RAND_3067 = {1{`RANDOM}};
  mesh_15_15_io_in_control_0_dataflow_pipe_b = _RAND_3067[0:0];
  _RAND_3068 = {1{`RANDOM}};
  mesh_15_15_io_in_control_0_propagate_pipe_b = _RAND_3068[0:0];
  _RAND_3069 = {1{`RANDOM}};
  mesh_15_15_io_in_control_1_shift_pipe_b = _RAND_3069[4:0];
  _RAND_3070 = {1{`RANDOM}};
  mesh_15_15_io_in_control_1_dataflow_pipe_b = _RAND_3070[0:0];
  _RAND_3071 = {1{`RANDOM}};
  mesh_15_15_io_in_control_1_propagate_pipe_b = _RAND_3071[0:0];
  _RAND_3072 = {1{`RANDOM}};
  r_256_0 = _RAND_3072[0:0];
  _RAND_3073 = {1{`RANDOM}};
  r_256_1 = _RAND_3073[0:0];
  _RAND_3074 = {1{`RANDOM}};
  r_257_0 = _RAND_3074[0:0];
  _RAND_3075 = {1{`RANDOM}};
  r_257_1 = _RAND_3075[0:0];
  _RAND_3076 = {1{`RANDOM}};
  r_258_0 = _RAND_3076[0:0];
  _RAND_3077 = {1{`RANDOM}};
  r_258_1 = _RAND_3077[0:0];
  _RAND_3078 = {1{`RANDOM}};
  r_259_0 = _RAND_3078[0:0];
  _RAND_3079 = {1{`RANDOM}};
  r_259_1 = _RAND_3079[0:0];
  _RAND_3080 = {1{`RANDOM}};
  r_260_0 = _RAND_3080[0:0];
  _RAND_3081 = {1{`RANDOM}};
  r_260_1 = _RAND_3081[0:0];
  _RAND_3082 = {1{`RANDOM}};
  r_261_0 = _RAND_3082[0:0];
  _RAND_3083 = {1{`RANDOM}};
  r_261_1 = _RAND_3083[0:0];
  _RAND_3084 = {1{`RANDOM}};
  r_262_0 = _RAND_3084[0:0];
  _RAND_3085 = {1{`RANDOM}};
  r_262_1 = _RAND_3085[0:0];
  _RAND_3086 = {1{`RANDOM}};
  r_263_0 = _RAND_3086[0:0];
  _RAND_3087 = {1{`RANDOM}};
  r_263_1 = _RAND_3087[0:0];
  _RAND_3088 = {1{`RANDOM}};
  r_264_0 = _RAND_3088[0:0];
  _RAND_3089 = {1{`RANDOM}};
  r_264_1 = _RAND_3089[0:0];
  _RAND_3090 = {1{`RANDOM}};
  r_265_0 = _RAND_3090[0:0];
  _RAND_3091 = {1{`RANDOM}};
  r_265_1 = _RAND_3091[0:0];
  _RAND_3092 = {1{`RANDOM}};
  r_266_0 = _RAND_3092[0:0];
  _RAND_3093 = {1{`RANDOM}};
  r_266_1 = _RAND_3093[0:0];
  _RAND_3094 = {1{`RANDOM}};
  r_267_0 = _RAND_3094[0:0];
  _RAND_3095 = {1{`RANDOM}};
  r_267_1 = _RAND_3095[0:0];
  _RAND_3096 = {1{`RANDOM}};
  r_268_0 = _RAND_3096[0:0];
  _RAND_3097 = {1{`RANDOM}};
  r_268_1 = _RAND_3097[0:0];
  _RAND_3098 = {1{`RANDOM}};
  r_269_0 = _RAND_3098[0:0];
  _RAND_3099 = {1{`RANDOM}};
  r_269_1 = _RAND_3099[0:0];
  _RAND_3100 = {1{`RANDOM}};
  r_270_0 = _RAND_3100[0:0];
  _RAND_3101 = {1{`RANDOM}};
  r_270_1 = _RAND_3101[0:0];
  _RAND_3102 = {1{`RANDOM}};
  r_271_0 = _RAND_3102[0:0];
  _RAND_3103 = {1{`RANDOM}};
  r_271_1 = _RAND_3103[0:0];
  _RAND_3104 = {1{`RANDOM}};
  r_272_0 = _RAND_3104[0:0];
  _RAND_3105 = {1{`RANDOM}};
  r_272_1 = _RAND_3105[0:0];
  _RAND_3106 = {1{`RANDOM}};
  r_273_0 = _RAND_3106[0:0];
  _RAND_3107 = {1{`RANDOM}};
  r_273_1 = _RAND_3107[0:0];
  _RAND_3108 = {1{`RANDOM}};
  r_274_0 = _RAND_3108[0:0];
  _RAND_3109 = {1{`RANDOM}};
  r_274_1 = _RAND_3109[0:0];
  _RAND_3110 = {1{`RANDOM}};
  r_275_0 = _RAND_3110[0:0];
  _RAND_3111 = {1{`RANDOM}};
  r_275_1 = _RAND_3111[0:0];
  _RAND_3112 = {1{`RANDOM}};
  r_276_0 = _RAND_3112[0:0];
  _RAND_3113 = {1{`RANDOM}};
  r_276_1 = _RAND_3113[0:0];
  _RAND_3114 = {1{`RANDOM}};
  r_277_0 = _RAND_3114[0:0];
  _RAND_3115 = {1{`RANDOM}};
  r_277_1 = _RAND_3115[0:0];
  _RAND_3116 = {1{`RANDOM}};
  r_278_0 = _RAND_3116[0:0];
  _RAND_3117 = {1{`RANDOM}};
  r_278_1 = _RAND_3117[0:0];
  _RAND_3118 = {1{`RANDOM}};
  r_279_0 = _RAND_3118[0:0];
  _RAND_3119 = {1{`RANDOM}};
  r_279_1 = _RAND_3119[0:0];
  _RAND_3120 = {1{`RANDOM}};
  r_280_0 = _RAND_3120[0:0];
  _RAND_3121 = {1{`RANDOM}};
  r_280_1 = _RAND_3121[0:0];
  _RAND_3122 = {1{`RANDOM}};
  r_281_0 = _RAND_3122[0:0];
  _RAND_3123 = {1{`RANDOM}};
  r_281_1 = _RAND_3123[0:0];
  _RAND_3124 = {1{`RANDOM}};
  r_282_0 = _RAND_3124[0:0];
  _RAND_3125 = {1{`RANDOM}};
  r_282_1 = _RAND_3125[0:0];
  _RAND_3126 = {1{`RANDOM}};
  r_283_0 = _RAND_3126[0:0];
  _RAND_3127 = {1{`RANDOM}};
  r_283_1 = _RAND_3127[0:0];
  _RAND_3128 = {1{`RANDOM}};
  r_284_0 = _RAND_3128[0:0];
  _RAND_3129 = {1{`RANDOM}};
  r_284_1 = _RAND_3129[0:0];
  _RAND_3130 = {1{`RANDOM}};
  r_285_0 = _RAND_3130[0:0];
  _RAND_3131 = {1{`RANDOM}};
  r_285_1 = _RAND_3131[0:0];
  _RAND_3132 = {1{`RANDOM}};
  r_286_0 = _RAND_3132[0:0];
  _RAND_3133 = {1{`RANDOM}};
  r_286_1 = _RAND_3133[0:0];
  _RAND_3134 = {1{`RANDOM}};
  r_287_0 = _RAND_3134[0:0];
  _RAND_3135 = {1{`RANDOM}};
  r_287_1 = _RAND_3135[0:0];
  _RAND_3136 = {1{`RANDOM}};
  r_288_0 = _RAND_3136[0:0];
  _RAND_3137 = {1{`RANDOM}};
  r_288_1 = _RAND_3137[0:0];
  _RAND_3138 = {1{`RANDOM}};
  r_289_0 = _RAND_3138[0:0];
  _RAND_3139 = {1{`RANDOM}};
  r_289_1 = _RAND_3139[0:0];
  _RAND_3140 = {1{`RANDOM}};
  r_290_0 = _RAND_3140[0:0];
  _RAND_3141 = {1{`RANDOM}};
  r_290_1 = _RAND_3141[0:0];
  _RAND_3142 = {1{`RANDOM}};
  r_291_0 = _RAND_3142[0:0];
  _RAND_3143 = {1{`RANDOM}};
  r_291_1 = _RAND_3143[0:0];
  _RAND_3144 = {1{`RANDOM}};
  r_292_0 = _RAND_3144[0:0];
  _RAND_3145 = {1{`RANDOM}};
  r_292_1 = _RAND_3145[0:0];
  _RAND_3146 = {1{`RANDOM}};
  r_293_0 = _RAND_3146[0:0];
  _RAND_3147 = {1{`RANDOM}};
  r_293_1 = _RAND_3147[0:0];
  _RAND_3148 = {1{`RANDOM}};
  r_294_0 = _RAND_3148[0:0];
  _RAND_3149 = {1{`RANDOM}};
  r_294_1 = _RAND_3149[0:0];
  _RAND_3150 = {1{`RANDOM}};
  r_295_0 = _RAND_3150[0:0];
  _RAND_3151 = {1{`RANDOM}};
  r_295_1 = _RAND_3151[0:0];
  _RAND_3152 = {1{`RANDOM}};
  r_296_0 = _RAND_3152[0:0];
  _RAND_3153 = {1{`RANDOM}};
  r_296_1 = _RAND_3153[0:0];
  _RAND_3154 = {1{`RANDOM}};
  r_297_0 = _RAND_3154[0:0];
  _RAND_3155 = {1{`RANDOM}};
  r_297_1 = _RAND_3155[0:0];
  _RAND_3156 = {1{`RANDOM}};
  r_298_0 = _RAND_3156[0:0];
  _RAND_3157 = {1{`RANDOM}};
  r_298_1 = _RAND_3157[0:0];
  _RAND_3158 = {1{`RANDOM}};
  r_299_0 = _RAND_3158[0:0];
  _RAND_3159 = {1{`RANDOM}};
  r_299_1 = _RAND_3159[0:0];
  _RAND_3160 = {1{`RANDOM}};
  r_300_0 = _RAND_3160[0:0];
  _RAND_3161 = {1{`RANDOM}};
  r_300_1 = _RAND_3161[0:0];
  _RAND_3162 = {1{`RANDOM}};
  r_301_0 = _RAND_3162[0:0];
  _RAND_3163 = {1{`RANDOM}};
  r_301_1 = _RAND_3163[0:0];
  _RAND_3164 = {1{`RANDOM}};
  r_302_0 = _RAND_3164[0:0];
  _RAND_3165 = {1{`RANDOM}};
  r_302_1 = _RAND_3165[0:0];
  _RAND_3166 = {1{`RANDOM}};
  r_303_0 = _RAND_3166[0:0];
  _RAND_3167 = {1{`RANDOM}};
  r_303_1 = _RAND_3167[0:0];
  _RAND_3168 = {1{`RANDOM}};
  r_304_0 = _RAND_3168[0:0];
  _RAND_3169 = {1{`RANDOM}};
  r_304_1 = _RAND_3169[0:0];
  _RAND_3170 = {1{`RANDOM}};
  r_305_0 = _RAND_3170[0:0];
  _RAND_3171 = {1{`RANDOM}};
  r_305_1 = _RAND_3171[0:0];
  _RAND_3172 = {1{`RANDOM}};
  r_306_0 = _RAND_3172[0:0];
  _RAND_3173 = {1{`RANDOM}};
  r_306_1 = _RAND_3173[0:0];
  _RAND_3174 = {1{`RANDOM}};
  r_307_0 = _RAND_3174[0:0];
  _RAND_3175 = {1{`RANDOM}};
  r_307_1 = _RAND_3175[0:0];
  _RAND_3176 = {1{`RANDOM}};
  r_308_0 = _RAND_3176[0:0];
  _RAND_3177 = {1{`RANDOM}};
  r_308_1 = _RAND_3177[0:0];
  _RAND_3178 = {1{`RANDOM}};
  r_309_0 = _RAND_3178[0:0];
  _RAND_3179 = {1{`RANDOM}};
  r_309_1 = _RAND_3179[0:0];
  _RAND_3180 = {1{`RANDOM}};
  r_310_0 = _RAND_3180[0:0];
  _RAND_3181 = {1{`RANDOM}};
  r_310_1 = _RAND_3181[0:0];
  _RAND_3182 = {1{`RANDOM}};
  r_311_0 = _RAND_3182[0:0];
  _RAND_3183 = {1{`RANDOM}};
  r_311_1 = _RAND_3183[0:0];
  _RAND_3184 = {1{`RANDOM}};
  r_312_0 = _RAND_3184[0:0];
  _RAND_3185 = {1{`RANDOM}};
  r_312_1 = _RAND_3185[0:0];
  _RAND_3186 = {1{`RANDOM}};
  r_313_0 = _RAND_3186[0:0];
  _RAND_3187 = {1{`RANDOM}};
  r_313_1 = _RAND_3187[0:0];
  _RAND_3188 = {1{`RANDOM}};
  r_314_0 = _RAND_3188[0:0];
  _RAND_3189 = {1{`RANDOM}};
  r_314_1 = _RAND_3189[0:0];
  _RAND_3190 = {1{`RANDOM}};
  r_315_0 = _RAND_3190[0:0];
  _RAND_3191 = {1{`RANDOM}};
  r_315_1 = _RAND_3191[0:0];
  _RAND_3192 = {1{`RANDOM}};
  r_316_0 = _RAND_3192[0:0];
  _RAND_3193 = {1{`RANDOM}};
  r_316_1 = _RAND_3193[0:0];
  _RAND_3194 = {1{`RANDOM}};
  r_317_0 = _RAND_3194[0:0];
  _RAND_3195 = {1{`RANDOM}};
  r_317_1 = _RAND_3195[0:0];
  _RAND_3196 = {1{`RANDOM}};
  r_318_0 = _RAND_3196[0:0];
  _RAND_3197 = {1{`RANDOM}};
  r_318_1 = _RAND_3197[0:0];
  _RAND_3198 = {1{`RANDOM}};
  r_319_0 = _RAND_3198[0:0];
  _RAND_3199 = {1{`RANDOM}};
  r_319_1 = _RAND_3199[0:0];
  _RAND_3200 = {1{`RANDOM}};
  r_320_0 = _RAND_3200[0:0];
  _RAND_3201 = {1{`RANDOM}};
  r_320_1 = _RAND_3201[0:0];
  _RAND_3202 = {1{`RANDOM}};
  r_321_0 = _RAND_3202[0:0];
  _RAND_3203 = {1{`RANDOM}};
  r_321_1 = _RAND_3203[0:0];
  _RAND_3204 = {1{`RANDOM}};
  r_322_0 = _RAND_3204[0:0];
  _RAND_3205 = {1{`RANDOM}};
  r_322_1 = _RAND_3205[0:0];
  _RAND_3206 = {1{`RANDOM}};
  r_323_0 = _RAND_3206[0:0];
  _RAND_3207 = {1{`RANDOM}};
  r_323_1 = _RAND_3207[0:0];
  _RAND_3208 = {1{`RANDOM}};
  r_324_0 = _RAND_3208[0:0];
  _RAND_3209 = {1{`RANDOM}};
  r_324_1 = _RAND_3209[0:0];
  _RAND_3210 = {1{`RANDOM}};
  r_325_0 = _RAND_3210[0:0];
  _RAND_3211 = {1{`RANDOM}};
  r_325_1 = _RAND_3211[0:0];
  _RAND_3212 = {1{`RANDOM}};
  r_326_0 = _RAND_3212[0:0];
  _RAND_3213 = {1{`RANDOM}};
  r_326_1 = _RAND_3213[0:0];
  _RAND_3214 = {1{`RANDOM}};
  r_327_0 = _RAND_3214[0:0];
  _RAND_3215 = {1{`RANDOM}};
  r_327_1 = _RAND_3215[0:0];
  _RAND_3216 = {1{`RANDOM}};
  r_328_0 = _RAND_3216[0:0];
  _RAND_3217 = {1{`RANDOM}};
  r_328_1 = _RAND_3217[0:0];
  _RAND_3218 = {1{`RANDOM}};
  r_329_0 = _RAND_3218[0:0];
  _RAND_3219 = {1{`RANDOM}};
  r_329_1 = _RAND_3219[0:0];
  _RAND_3220 = {1{`RANDOM}};
  r_330_0 = _RAND_3220[0:0];
  _RAND_3221 = {1{`RANDOM}};
  r_330_1 = _RAND_3221[0:0];
  _RAND_3222 = {1{`RANDOM}};
  r_331_0 = _RAND_3222[0:0];
  _RAND_3223 = {1{`RANDOM}};
  r_331_1 = _RAND_3223[0:0];
  _RAND_3224 = {1{`RANDOM}};
  r_332_0 = _RAND_3224[0:0];
  _RAND_3225 = {1{`RANDOM}};
  r_332_1 = _RAND_3225[0:0];
  _RAND_3226 = {1{`RANDOM}};
  r_333_0 = _RAND_3226[0:0];
  _RAND_3227 = {1{`RANDOM}};
  r_333_1 = _RAND_3227[0:0];
  _RAND_3228 = {1{`RANDOM}};
  r_334_0 = _RAND_3228[0:0];
  _RAND_3229 = {1{`RANDOM}};
  r_334_1 = _RAND_3229[0:0];
  _RAND_3230 = {1{`RANDOM}};
  r_335_0 = _RAND_3230[0:0];
  _RAND_3231 = {1{`RANDOM}};
  r_335_1 = _RAND_3231[0:0];
  _RAND_3232 = {1{`RANDOM}};
  r_336_0 = _RAND_3232[0:0];
  _RAND_3233 = {1{`RANDOM}};
  r_336_1 = _RAND_3233[0:0];
  _RAND_3234 = {1{`RANDOM}};
  r_337_0 = _RAND_3234[0:0];
  _RAND_3235 = {1{`RANDOM}};
  r_337_1 = _RAND_3235[0:0];
  _RAND_3236 = {1{`RANDOM}};
  r_338_0 = _RAND_3236[0:0];
  _RAND_3237 = {1{`RANDOM}};
  r_338_1 = _RAND_3237[0:0];
  _RAND_3238 = {1{`RANDOM}};
  r_339_0 = _RAND_3238[0:0];
  _RAND_3239 = {1{`RANDOM}};
  r_339_1 = _RAND_3239[0:0];
  _RAND_3240 = {1{`RANDOM}};
  r_340_0 = _RAND_3240[0:0];
  _RAND_3241 = {1{`RANDOM}};
  r_340_1 = _RAND_3241[0:0];
  _RAND_3242 = {1{`RANDOM}};
  r_341_0 = _RAND_3242[0:0];
  _RAND_3243 = {1{`RANDOM}};
  r_341_1 = _RAND_3243[0:0];
  _RAND_3244 = {1{`RANDOM}};
  r_342_0 = _RAND_3244[0:0];
  _RAND_3245 = {1{`RANDOM}};
  r_342_1 = _RAND_3245[0:0];
  _RAND_3246 = {1{`RANDOM}};
  r_343_0 = _RAND_3246[0:0];
  _RAND_3247 = {1{`RANDOM}};
  r_343_1 = _RAND_3247[0:0];
  _RAND_3248 = {1{`RANDOM}};
  r_344_0 = _RAND_3248[0:0];
  _RAND_3249 = {1{`RANDOM}};
  r_344_1 = _RAND_3249[0:0];
  _RAND_3250 = {1{`RANDOM}};
  r_345_0 = _RAND_3250[0:0];
  _RAND_3251 = {1{`RANDOM}};
  r_345_1 = _RAND_3251[0:0];
  _RAND_3252 = {1{`RANDOM}};
  r_346_0 = _RAND_3252[0:0];
  _RAND_3253 = {1{`RANDOM}};
  r_346_1 = _RAND_3253[0:0];
  _RAND_3254 = {1{`RANDOM}};
  r_347_0 = _RAND_3254[0:0];
  _RAND_3255 = {1{`RANDOM}};
  r_347_1 = _RAND_3255[0:0];
  _RAND_3256 = {1{`RANDOM}};
  r_348_0 = _RAND_3256[0:0];
  _RAND_3257 = {1{`RANDOM}};
  r_348_1 = _RAND_3257[0:0];
  _RAND_3258 = {1{`RANDOM}};
  r_349_0 = _RAND_3258[0:0];
  _RAND_3259 = {1{`RANDOM}};
  r_349_1 = _RAND_3259[0:0];
  _RAND_3260 = {1{`RANDOM}};
  r_350_0 = _RAND_3260[0:0];
  _RAND_3261 = {1{`RANDOM}};
  r_350_1 = _RAND_3261[0:0];
  _RAND_3262 = {1{`RANDOM}};
  r_351_0 = _RAND_3262[0:0];
  _RAND_3263 = {1{`RANDOM}};
  r_351_1 = _RAND_3263[0:0];
  _RAND_3264 = {1{`RANDOM}};
  r_352_0 = _RAND_3264[0:0];
  _RAND_3265 = {1{`RANDOM}};
  r_352_1 = _RAND_3265[0:0];
  _RAND_3266 = {1{`RANDOM}};
  r_353_0 = _RAND_3266[0:0];
  _RAND_3267 = {1{`RANDOM}};
  r_353_1 = _RAND_3267[0:0];
  _RAND_3268 = {1{`RANDOM}};
  r_354_0 = _RAND_3268[0:0];
  _RAND_3269 = {1{`RANDOM}};
  r_354_1 = _RAND_3269[0:0];
  _RAND_3270 = {1{`RANDOM}};
  r_355_0 = _RAND_3270[0:0];
  _RAND_3271 = {1{`RANDOM}};
  r_355_1 = _RAND_3271[0:0];
  _RAND_3272 = {1{`RANDOM}};
  r_356_0 = _RAND_3272[0:0];
  _RAND_3273 = {1{`RANDOM}};
  r_356_1 = _RAND_3273[0:0];
  _RAND_3274 = {1{`RANDOM}};
  r_357_0 = _RAND_3274[0:0];
  _RAND_3275 = {1{`RANDOM}};
  r_357_1 = _RAND_3275[0:0];
  _RAND_3276 = {1{`RANDOM}};
  r_358_0 = _RAND_3276[0:0];
  _RAND_3277 = {1{`RANDOM}};
  r_358_1 = _RAND_3277[0:0];
  _RAND_3278 = {1{`RANDOM}};
  r_359_0 = _RAND_3278[0:0];
  _RAND_3279 = {1{`RANDOM}};
  r_359_1 = _RAND_3279[0:0];
  _RAND_3280 = {1{`RANDOM}};
  r_360_0 = _RAND_3280[0:0];
  _RAND_3281 = {1{`RANDOM}};
  r_360_1 = _RAND_3281[0:0];
  _RAND_3282 = {1{`RANDOM}};
  r_361_0 = _RAND_3282[0:0];
  _RAND_3283 = {1{`RANDOM}};
  r_361_1 = _RAND_3283[0:0];
  _RAND_3284 = {1{`RANDOM}};
  r_362_0 = _RAND_3284[0:0];
  _RAND_3285 = {1{`RANDOM}};
  r_362_1 = _RAND_3285[0:0];
  _RAND_3286 = {1{`RANDOM}};
  r_363_0 = _RAND_3286[0:0];
  _RAND_3287 = {1{`RANDOM}};
  r_363_1 = _RAND_3287[0:0];
  _RAND_3288 = {1{`RANDOM}};
  r_364_0 = _RAND_3288[0:0];
  _RAND_3289 = {1{`RANDOM}};
  r_364_1 = _RAND_3289[0:0];
  _RAND_3290 = {1{`RANDOM}};
  r_365_0 = _RAND_3290[0:0];
  _RAND_3291 = {1{`RANDOM}};
  r_365_1 = _RAND_3291[0:0];
  _RAND_3292 = {1{`RANDOM}};
  r_366_0 = _RAND_3292[0:0];
  _RAND_3293 = {1{`RANDOM}};
  r_366_1 = _RAND_3293[0:0];
  _RAND_3294 = {1{`RANDOM}};
  r_367_0 = _RAND_3294[0:0];
  _RAND_3295 = {1{`RANDOM}};
  r_367_1 = _RAND_3295[0:0];
  _RAND_3296 = {1{`RANDOM}};
  r_368_0 = _RAND_3296[0:0];
  _RAND_3297 = {1{`RANDOM}};
  r_368_1 = _RAND_3297[0:0];
  _RAND_3298 = {1{`RANDOM}};
  r_369_0 = _RAND_3298[0:0];
  _RAND_3299 = {1{`RANDOM}};
  r_369_1 = _RAND_3299[0:0];
  _RAND_3300 = {1{`RANDOM}};
  r_370_0 = _RAND_3300[0:0];
  _RAND_3301 = {1{`RANDOM}};
  r_370_1 = _RAND_3301[0:0];
  _RAND_3302 = {1{`RANDOM}};
  r_371_0 = _RAND_3302[0:0];
  _RAND_3303 = {1{`RANDOM}};
  r_371_1 = _RAND_3303[0:0];
  _RAND_3304 = {1{`RANDOM}};
  r_372_0 = _RAND_3304[0:0];
  _RAND_3305 = {1{`RANDOM}};
  r_372_1 = _RAND_3305[0:0];
  _RAND_3306 = {1{`RANDOM}};
  r_373_0 = _RAND_3306[0:0];
  _RAND_3307 = {1{`RANDOM}};
  r_373_1 = _RAND_3307[0:0];
  _RAND_3308 = {1{`RANDOM}};
  r_374_0 = _RAND_3308[0:0];
  _RAND_3309 = {1{`RANDOM}};
  r_374_1 = _RAND_3309[0:0];
  _RAND_3310 = {1{`RANDOM}};
  r_375_0 = _RAND_3310[0:0];
  _RAND_3311 = {1{`RANDOM}};
  r_375_1 = _RAND_3311[0:0];
  _RAND_3312 = {1{`RANDOM}};
  r_376_0 = _RAND_3312[0:0];
  _RAND_3313 = {1{`RANDOM}};
  r_376_1 = _RAND_3313[0:0];
  _RAND_3314 = {1{`RANDOM}};
  r_377_0 = _RAND_3314[0:0];
  _RAND_3315 = {1{`RANDOM}};
  r_377_1 = _RAND_3315[0:0];
  _RAND_3316 = {1{`RANDOM}};
  r_378_0 = _RAND_3316[0:0];
  _RAND_3317 = {1{`RANDOM}};
  r_378_1 = _RAND_3317[0:0];
  _RAND_3318 = {1{`RANDOM}};
  r_379_0 = _RAND_3318[0:0];
  _RAND_3319 = {1{`RANDOM}};
  r_379_1 = _RAND_3319[0:0];
  _RAND_3320 = {1{`RANDOM}};
  r_380_0 = _RAND_3320[0:0];
  _RAND_3321 = {1{`RANDOM}};
  r_380_1 = _RAND_3321[0:0];
  _RAND_3322 = {1{`RANDOM}};
  r_381_0 = _RAND_3322[0:0];
  _RAND_3323 = {1{`RANDOM}};
  r_381_1 = _RAND_3323[0:0];
  _RAND_3324 = {1{`RANDOM}};
  r_382_0 = _RAND_3324[0:0];
  _RAND_3325 = {1{`RANDOM}};
  r_382_1 = _RAND_3325[0:0];
  _RAND_3326 = {1{`RANDOM}};
  r_383_0 = _RAND_3326[0:0];
  _RAND_3327 = {1{`RANDOM}};
  r_383_1 = _RAND_3327[0:0];
  _RAND_3328 = {1{`RANDOM}};
  r_384_0 = _RAND_3328[0:0];
  _RAND_3329 = {1{`RANDOM}};
  r_384_1 = _RAND_3329[0:0];
  _RAND_3330 = {1{`RANDOM}};
  r_385_0 = _RAND_3330[0:0];
  _RAND_3331 = {1{`RANDOM}};
  r_385_1 = _RAND_3331[0:0];
  _RAND_3332 = {1{`RANDOM}};
  r_386_0 = _RAND_3332[0:0];
  _RAND_3333 = {1{`RANDOM}};
  r_386_1 = _RAND_3333[0:0];
  _RAND_3334 = {1{`RANDOM}};
  r_387_0 = _RAND_3334[0:0];
  _RAND_3335 = {1{`RANDOM}};
  r_387_1 = _RAND_3335[0:0];
  _RAND_3336 = {1{`RANDOM}};
  r_388_0 = _RAND_3336[0:0];
  _RAND_3337 = {1{`RANDOM}};
  r_388_1 = _RAND_3337[0:0];
  _RAND_3338 = {1{`RANDOM}};
  r_389_0 = _RAND_3338[0:0];
  _RAND_3339 = {1{`RANDOM}};
  r_389_1 = _RAND_3339[0:0];
  _RAND_3340 = {1{`RANDOM}};
  r_390_0 = _RAND_3340[0:0];
  _RAND_3341 = {1{`RANDOM}};
  r_390_1 = _RAND_3341[0:0];
  _RAND_3342 = {1{`RANDOM}};
  r_391_0 = _RAND_3342[0:0];
  _RAND_3343 = {1{`RANDOM}};
  r_391_1 = _RAND_3343[0:0];
  _RAND_3344 = {1{`RANDOM}};
  r_392_0 = _RAND_3344[0:0];
  _RAND_3345 = {1{`RANDOM}};
  r_392_1 = _RAND_3345[0:0];
  _RAND_3346 = {1{`RANDOM}};
  r_393_0 = _RAND_3346[0:0];
  _RAND_3347 = {1{`RANDOM}};
  r_393_1 = _RAND_3347[0:0];
  _RAND_3348 = {1{`RANDOM}};
  r_394_0 = _RAND_3348[0:0];
  _RAND_3349 = {1{`RANDOM}};
  r_394_1 = _RAND_3349[0:0];
  _RAND_3350 = {1{`RANDOM}};
  r_395_0 = _RAND_3350[0:0];
  _RAND_3351 = {1{`RANDOM}};
  r_395_1 = _RAND_3351[0:0];
  _RAND_3352 = {1{`RANDOM}};
  r_396_0 = _RAND_3352[0:0];
  _RAND_3353 = {1{`RANDOM}};
  r_396_1 = _RAND_3353[0:0];
  _RAND_3354 = {1{`RANDOM}};
  r_397_0 = _RAND_3354[0:0];
  _RAND_3355 = {1{`RANDOM}};
  r_397_1 = _RAND_3355[0:0];
  _RAND_3356 = {1{`RANDOM}};
  r_398_0 = _RAND_3356[0:0];
  _RAND_3357 = {1{`RANDOM}};
  r_398_1 = _RAND_3357[0:0];
  _RAND_3358 = {1{`RANDOM}};
  r_399_0 = _RAND_3358[0:0];
  _RAND_3359 = {1{`RANDOM}};
  r_399_1 = _RAND_3359[0:0];
  _RAND_3360 = {1{`RANDOM}};
  r_400_0 = _RAND_3360[0:0];
  _RAND_3361 = {1{`RANDOM}};
  r_400_1 = _RAND_3361[0:0];
  _RAND_3362 = {1{`RANDOM}};
  r_401_0 = _RAND_3362[0:0];
  _RAND_3363 = {1{`RANDOM}};
  r_401_1 = _RAND_3363[0:0];
  _RAND_3364 = {1{`RANDOM}};
  r_402_0 = _RAND_3364[0:0];
  _RAND_3365 = {1{`RANDOM}};
  r_402_1 = _RAND_3365[0:0];
  _RAND_3366 = {1{`RANDOM}};
  r_403_0 = _RAND_3366[0:0];
  _RAND_3367 = {1{`RANDOM}};
  r_403_1 = _RAND_3367[0:0];
  _RAND_3368 = {1{`RANDOM}};
  r_404_0 = _RAND_3368[0:0];
  _RAND_3369 = {1{`RANDOM}};
  r_404_1 = _RAND_3369[0:0];
  _RAND_3370 = {1{`RANDOM}};
  r_405_0 = _RAND_3370[0:0];
  _RAND_3371 = {1{`RANDOM}};
  r_405_1 = _RAND_3371[0:0];
  _RAND_3372 = {1{`RANDOM}};
  r_406_0 = _RAND_3372[0:0];
  _RAND_3373 = {1{`RANDOM}};
  r_406_1 = _RAND_3373[0:0];
  _RAND_3374 = {1{`RANDOM}};
  r_407_0 = _RAND_3374[0:0];
  _RAND_3375 = {1{`RANDOM}};
  r_407_1 = _RAND_3375[0:0];
  _RAND_3376 = {1{`RANDOM}};
  r_408_0 = _RAND_3376[0:0];
  _RAND_3377 = {1{`RANDOM}};
  r_408_1 = _RAND_3377[0:0];
  _RAND_3378 = {1{`RANDOM}};
  r_409_0 = _RAND_3378[0:0];
  _RAND_3379 = {1{`RANDOM}};
  r_409_1 = _RAND_3379[0:0];
  _RAND_3380 = {1{`RANDOM}};
  r_410_0 = _RAND_3380[0:0];
  _RAND_3381 = {1{`RANDOM}};
  r_410_1 = _RAND_3381[0:0];
  _RAND_3382 = {1{`RANDOM}};
  r_411_0 = _RAND_3382[0:0];
  _RAND_3383 = {1{`RANDOM}};
  r_411_1 = _RAND_3383[0:0];
  _RAND_3384 = {1{`RANDOM}};
  r_412_0 = _RAND_3384[0:0];
  _RAND_3385 = {1{`RANDOM}};
  r_412_1 = _RAND_3385[0:0];
  _RAND_3386 = {1{`RANDOM}};
  r_413_0 = _RAND_3386[0:0];
  _RAND_3387 = {1{`RANDOM}};
  r_413_1 = _RAND_3387[0:0];
  _RAND_3388 = {1{`RANDOM}};
  r_414_0 = _RAND_3388[0:0];
  _RAND_3389 = {1{`RANDOM}};
  r_414_1 = _RAND_3389[0:0];
  _RAND_3390 = {1{`RANDOM}};
  r_415_0 = _RAND_3390[0:0];
  _RAND_3391 = {1{`RANDOM}};
  r_415_1 = _RAND_3391[0:0];
  _RAND_3392 = {1{`RANDOM}};
  r_416_0 = _RAND_3392[0:0];
  _RAND_3393 = {1{`RANDOM}};
  r_416_1 = _RAND_3393[0:0];
  _RAND_3394 = {1{`RANDOM}};
  r_417_0 = _RAND_3394[0:0];
  _RAND_3395 = {1{`RANDOM}};
  r_417_1 = _RAND_3395[0:0];
  _RAND_3396 = {1{`RANDOM}};
  r_418_0 = _RAND_3396[0:0];
  _RAND_3397 = {1{`RANDOM}};
  r_418_1 = _RAND_3397[0:0];
  _RAND_3398 = {1{`RANDOM}};
  r_419_0 = _RAND_3398[0:0];
  _RAND_3399 = {1{`RANDOM}};
  r_419_1 = _RAND_3399[0:0];
  _RAND_3400 = {1{`RANDOM}};
  r_420_0 = _RAND_3400[0:0];
  _RAND_3401 = {1{`RANDOM}};
  r_420_1 = _RAND_3401[0:0];
  _RAND_3402 = {1{`RANDOM}};
  r_421_0 = _RAND_3402[0:0];
  _RAND_3403 = {1{`RANDOM}};
  r_421_1 = _RAND_3403[0:0];
  _RAND_3404 = {1{`RANDOM}};
  r_422_0 = _RAND_3404[0:0];
  _RAND_3405 = {1{`RANDOM}};
  r_422_1 = _RAND_3405[0:0];
  _RAND_3406 = {1{`RANDOM}};
  r_423_0 = _RAND_3406[0:0];
  _RAND_3407 = {1{`RANDOM}};
  r_423_1 = _RAND_3407[0:0];
  _RAND_3408 = {1{`RANDOM}};
  r_424_0 = _RAND_3408[0:0];
  _RAND_3409 = {1{`RANDOM}};
  r_424_1 = _RAND_3409[0:0];
  _RAND_3410 = {1{`RANDOM}};
  r_425_0 = _RAND_3410[0:0];
  _RAND_3411 = {1{`RANDOM}};
  r_425_1 = _RAND_3411[0:0];
  _RAND_3412 = {1{`RANDOM}};
  r_426_0 = _RAND_3412[0:0];
  _RAND_3413 = {1{`RANDOM}};
  r_426_1 = _RAND_3413[0:0];
  _RAND_3414 = {1{`RANDOM}};
  r_427_0 = _RAND_3414[0:0];
  _RAND_3415 = {1{`RANDOM}};
  r_427_1 = _RAND_3415[0:0];
  _RAND_3416 = {1{`RANDOM}};
  r_428_0 = _RAND_3416[0:0];
  _RAND_3417 = {1{`RANDOM}};
  r_428_1 = _RAND_3417[0:0];
  _RAND_3418 = {1{`RANDOM}};
  r_429_0 = _RAND_3418[0:0];
  _RAND_3419 = {1{`RANDOM}};
  r_429_1 = _RAND_3419[0:0];
  _RAND_3420 = {1{`RANDOM}};
  r_430_0 = _RAND_3420[0:0];
  _RAND_3421 = {1{`RANDOM}};
  r_430_1 = _RAND_3421[0:0];
  _RAND_3422 = {1{`RANDOM}};
  r_431_0 = _RAND_3422[0:0];
  _RAND_3423 = {1{`RANDOM}};
  r_431_1 = _RAND_3423[0:0];
  _RAND_3424 = {1{`RANDOM}};
  r_432_0 = _RAND_3424[0:0];
  _RAND_3425 = {1{`RANDOM}};
  r_432_1 = _RAND_3425[0:0];
  _RAND_3426 = {1{`RANDOM}};
  r_433_0 = _RAND_3426[0:0];
  _RAND_3427 = {1{`RANDOM}};
  r_433_1 = _RAND_3427[0:0];
  _RAND_3428 = {1{`RANDOM}};
  r_434_0 = _RAND_3428[0:0];
  _RAND_3429 = {1{`RANDOM}};
  r_434_1 = _RAND_3429[0:0];
  _RAND_3430 = {1{`RANDOM}};
  r_435_0 = _RAND_3430[0:0];
  _RAND_3431 = {1{`RANDOM}};
  r_435_1 = _RAND_3431[0:0];
  _RAND_3432 = {1{`RANDOM}};
  r_436_0 = _RAND_3432[0:0];
  _RAND_3433 = {1{`RANDOM}};
  r_436_1 = _RAND_3433[0:0];
  _RAND_3434 = {1{`RANDOM}};
  r_437_0 = _RAND_3434[0:0];
  _RAND_3435 = {1{`RANDOM}};
  r_437_1 = _RAND_3435[0:0];
  _RAND_3436 = {1{`RANDOM}};
  r_438_0 = _RAND_3436[0:0];
  _RAND_3437 = {1{`RANDOM}};
  r_438_1 = _RAND_3437[0:0];
  _RAND_3438 = {1{`RANDOM}};
  r_439_0 = _RAND_3438[0:0];
  _RAND_3439 = {1{`RANDOM}};
  r_439_1 = _RAND_3439[0:0];
  _RAND_3440 = {1{`RANDOM}};
  r_440_0 = _RAND_3440[0:0];
  _RAND_3441 = {1{`RANDOM}};
  r_440_1 = _RAND_3441[0:0];
  _RAND_3442 = {1{`RANDOM}};
  r_441_0 = _RAND_3442[0:0];
  _RAND_3443 = {1{`RANDOM}};
  r_441_1 = _RAND_3443[0:0];
  _RAND_3444 = {1{`RANDOM}};
  r_442_0 = _RAND_3444[0:0];
  _RAND_3445 = {1{`RANDOM}};
  r_442_1 = _RAND_3445[0:0];
  _RAND_3446 = {1{`RANDOM}};
  r_443_0 = _RAND_3446[0:0];
  _RAND_3447 = {1{`RANDOM}};
  r_443_1 = _RAND_3447[0:0];
  _RAND_3448 = {1{`RANDOM}};
  r_444_0 = _RAND_3448[0:0];
  _RAND_3449 = {1{`RANDOM}};
  r_444_1 = _RAND_3449[0:0];
  _RAND_3450 = {1{`RANDOM}};
  r_445_0 = _RAND_3450[0:0];
  _RAND_3451 = {1{`RANDOM}};
  r_445_1 = _RAND_3451[0:0];
  _RAND_3452 = {1{`RANDOM}};
  r_446_0 = _RAND_3452[0:0];
  _RAND_3453 = {1{`RANDOM}};
  r_446_1 = _RAND_3453[0:0];
  _RAND_3454 = {1{`RANDOM}};
  r_447_0 = _RAND_3454[0:0];
  _RAND_3455 = {1{`RANDOM}};
  r_447_1 = _RAND_3455[0:0];
  _RAND_3456 = {1{`RANDOM}};
  r_448_0 = _RAND_3456[0:0];
  _RAND_3457 = {1{`RANDOM}};
  r_448_1 = _RAND_3457[0:0];
  _RAND_3458 = {1{`RANDOM}};
  r_449_0 = _RAND_3458[0:0];
  _RAND_3459 = {1{`RANDOM}};
  r_449_1 = _RAND_3459[0:0];
  _RAND_3460 = {1{`RANDOM}};
  r_450_0 = _RAND_3460[0:0];
  _RAND_3461 = {1{`RANDOM}};
  r_450_1 = _RAND_3461[0:0];
  _RAND_3462 = {1{`RANDOM}};
  r_451_0 = _RAND_3462[0:0];
  _RAND_3463 = {1{`RANDOM}};
  r_451_1 = _RAND_3463[0:0];
  _RAND_3464 = {1{`RANDOM}};
  r_452_0 = _RAND_3464[0:0];
  _RAND_3465 = {1{`RANDOM}};
  r_452_1 = _RAND_3465[0:0];
  _RAND_3466 = {1{`RANDOM}};
  r_453_0 = _RAND_3466[0:0];
  _RAND_3467 = {1{`RANDOM}};
  r_453_1 = _RAND_3467[0:0];
  _RAND_3468 = {1{`RANDOM}};
  r_454_0 = _RAND_3468[0:0];
  _RAND_3469 = {1{`RANDOM}};
  r_454_1 = _RAND_3469[0:0];
  _RAND_3470 = {1{`RANDOM}};
  r_455_0 = _RAND_3470[0:0];
  _RAND_3471 = {1{`RANDOM}};
  r_455_1 = _RAND_3471[0:0];
  _RAND_3472 = {1{`RANDOM}};
  r_456_0 = _RAND_3472[0:0];
  _RAND_3473 = {1{`RANDOM}};
  r_456_1 = _RAND_3473[0:0];
  _RAND_3474 = {1{`RANDOM}};
  r_457_0 = _RAND_3474[0:0];
  _RAND_3475 = {1{`RANDOM}};
  r_457_1 = _RAND_3475[0:0];
  _RAND_3476 = {1{`RANDOM}};
  r_458_0 = _RAND_3476[0:0];
  _RAND_3477 = {1{`RANDOM}};
  r_458_1 = _RAND_3477[0:0];
  _RAND_3478 = {1{`RANDOM}};
  r_459_0 = _RAND_3478[0:0];
  _RAND_3479 = {1{`RANDOM}};
  r_459_1 = _RAND_3479[0:0];
  _RAND_3480 = {1{`RANDOM}};
  r_460_0 = _RAND_3480[0:0];
  _RAND_3481 = {1{`RANDOM}};
  r_460_1 = _RAND_3481[0:0];
  _RAND_3482 = {1{`RANDOM}};
  r_461_0 = _RAND_3482[0:0];
  _RAND_3483 = {1{`RANDOM}};
  r_461_1 = _RAND_3483[0:0];
  _RAND_3484 = {1{`RANDOM}};
  r_462_0 = _RAND_3484[0:0];
  _RAND_3485 = {1{`RANDOM}};
  r_462_1 = _RAND_3485[0:0];
  _RAND_3486 = {1{`RANDOM}};
  r_463_0 = _RAND_3486[0:0];
  _RAND_3487 = {1{`RANDOM}};
  r_463_1 = _RAND_3487[0:0];
  _RAND_3488 = {1{`RANDOM}};
  r_464_0 = _RAND_3488[0:0];
  _RAND_3489 = {1{`RANDOM}};
  r_464_1 = _RAND_3489[0:0];
  _RAND_3490 = {1{`RANDOM}};
  r_465_0 = _RAND_3490[0:0];
  _RAND_3491 = {1{`RANDOM}};
  r_465_1 = _RAND_3491[0:0];
  _RAND_3492 = {1{`RANDOM}};
  r_466_0 = _RAND_3492[0:0];
  _RAND_3493 = {1{`RANDOM}};
  r_466_1 = _RAND_3493[0:0];
  _RAND_3494 = {1{`RANDOM}};
  r_467_0 = _RAND_3494[0:0];
  _RAND_3495 = {1{`RANDOM}};
  r_467_1 = _RAND_3495[0:0];
  _RAND_3496 = {1{`RANDOM}};
  r_468_0 = _RAND_3496[0:0];
  _RAND_3497 = {1{`RANDOM}};
  r_468_1 = _RAND_3497[0:0];
  _RAND_3498 = {1{`RANDOM}};
  r_469_0 = _RAND_3498[0:0];
  _RAND_3499 = {1{`RANDOM}};
  r_469_1 = _RAND_3499[0:0];
  _RAND_3500 = {1{`RANDOM}};
  r_470_0 = _RAND_3500[0:0];
  _RAND_3501 = {1{`RANDOM}};
  r_470_1 = _RAND_3501[0:0];
  _RAND_3502 = {1{`RANDOM}};
  r_471_0 = _RAND_3502[0:0];
  _RAND_3503 = {1{`RANDOM}};
  r_471_1 = _RAND_3503[0:0];
  _RAND_3504 = {1{`RANDOM}};
  r_472_0 = _RAND_3504[0:0];
  _RAND_3505 = {1{`RANDOM}};
  r_472_1 = _RAND_3505[0:0];
  _RAND_3506 = {1{`RANDOM}};
  r_473_0 = _RAND_3506[0:0];
  _RAND_3507 = {1{`RANDOM}};
  r_473_1 = _RAND_3507[0:0];
  _RAND_3508 = {1{`RANDOM}};
  r_474_0 = _RAND_3508[0:0];
  _RAND_3509 = {1{`RANDOM}};
  r_474_1 = _RAND_3509[0:0];
  _RAND_3510 = {1{`RANDOM}};
  r_475_0 = _RAND_3510[0:0];
  _RAND_3511 = {1{`RANDOM}};
  r_475_1 = _RAND_3511[0:0];
  _RAND_3512 = {1{`RANDOM}};
  r_476_0 = _RAND_3512[0:0];
  _RAND_3513 = {1{`RANDOM}};
  r_476_1 = _RAND_3513[0:0];
  _RAND_3514 = {1{`RANDOM}};
  r_477_0 = _RAND_3514[0:0];
  _RAND_3515 = {1{`RANDOM}};
  r_477_1 = _RAND_3515[0:0];
  _RAND_3516 = {1{`RANDOM}};
  r_478_0 = _RAND_3516[0:0];
  _RAND_3517 = {1{`RANDOM}};
  r_478_1 = _RAND_3517[0:0];
  _RAND_3518 = {1{`RANDOM}};
  r_479_0 = _RAND_3518[0:0];
  _RAND_3519 = {1{`RANDOM}};
  r_479_1 = _RAND_3519[0:0];
  _RAND_3520 = {1{`RANDOM}};
  r_480_0 = _RAND_3520[0:0];
  _RAND_3521 = {1{`RANDOM}};
  r_480_1 = _RAND_3521[0:0];
  _RAND_3522 = {1{`RANDOM}};
  r_481_0 = _RAND_3522[0:0];
  _RAND_3523 = {1{`RANDOM}};
  r_481_1 = _RAND_3523[0:0];
  _RAND_3524 = {1{`RANDOM}};
  r_482_0 = _RAND_3524[0:0];
  _RAND_3525 = {1{`RANDOM}};
  r_482_1 = _RAND_3525[0:0];
  _RAND_3526 = {1{`RANDOM}};
  r_483_0 = _RAND_3526[0:0];
  _RAND_3527 = {1{`RANDOM}};
  r_483_1 = _RAND_3527[0:0];
  _RAND_3528 = {1{`RANDOM}};
  r_484_0 = _RAND_3528[0:0];
  _RAND_3529 = {1{`RANDOM}};
  r_484_1 = _RAND_3529[0:0];
  _RAND_3530 = {1{`RANDOM}};
  r_485_0 = _RAND_3530[0:0];
  _RAND_3531 = {1{`RANDOM}};
  r_485_1 = _RAND_3531[0:0];
  _RAND_3532 = {1{`RANDOM}};
  r_486_0 = _RAND_3532[0:0];
  _RAND_3533 = {1{`RANDOM}};
  r_486_1 = _RAND_3533[0:0];
  _RAND_3534 = {1{`RANDOM}};
  r_487_0 = _RAND_3534[0:0];
  _RAND_3535 = {1{`RANDOM}};
  r_487_1 = _RAND_3535[0:0];
  _RAND_3536 = {1{`RANDOM}};
  r_488_0 = _RAND_3536[0:0];
  _RAND_3537 = {1{`RANDOM}};
  r_488_1 = _RAND_3537[0:0];
  _RAND_3538 = {1{`RANDOM}};
  r_489_0 = _RAND_3538[0:0];
  _RAND_3539 = {1{`RANDOM}};
  r_489_1 = _RAND_3539[0:0];
  _RAND_3540 = {1{`RANDOM}};
  r_490_0 = _RAND_3540[0:0];
  _RAND_3541 = {1{`RANDOM}};
  r_490_1 = _RAND_3541[0:0];
  _RAND_3542 = {1{`RANDOM}};
  r_491_0 = _RAND_3542[0:0];
  _RAND_3543 = {1{`RANDOM}};
  r_491_1 = _RAND_3543[0:0];
  _RAND_3544 = {1{`RANDOM}};
  r_492_0 = _RAND_3544[0:0];
  _RAND_3545 = {1{`RANDOM}};
  r_492_1 = _RAND_3545[0:0];
  _RAND_3546 = {1{`RANDOM}};
  r_493_0 = _RAND_3546[0:0];
  _RAND_3547 = {1{`RANDOM}};
  r_493_1 = _RAND_3547[0:0];
  _RAND_3548 = {1{`RANDOM}};
  r_494_0 = _RAND_3548[0:0];
  _RAND_3549 = {1{`RANDOM}};
  r_494_1 = _RAND_3549[0:0];
  _RAND_3550 = {1{`RANDOM}};
  r_495_0 = _RAND_3550[0:0];
  _RAND_3551 = {1{`RANDOM}};
  r_495_1 = _RAND_3551[0:0];
  _RAND_3552 = {1{`RANDOM}};
  r_496_0 = _RAND_3552[0:0];
  _RAND_3553 = {1{`RANDOM}};
  r_496_1 = _RAND_3553[0:0];
  _RAND_3554 = {1{`RANDOM}};
  r_497_0 = _RAND_3554[0:0];
  _RAND_3555 = {1{`RANDOM}};
  r_497_1 = _RAND_3555[0:0];
  _RAND_3556 = {1{`RANDOM}};
  r_498_0 = _RAND_3556[0:0];
  _RAND_3557 = {1{`RANDOM}};
  r_498_1 = _RAND_3557[0:0];
  _RAND_3558 = {1{`RANDOM}};
  r_499_0 = _RAND_3558[0:0];
  _RAND_3559 = {1{`RANDOM}};
  r_499_1 = _RAND_3559[0:0];
  _RAND_3560 = {1{`RANDOM}};
  r_500_0 = _RAND_3560[0:0];
  _RAND_3561 = {1{`RANDOM}};
  r_500_1 = _RAND_3561[0:0];
  _RAND_3562 = {1{`RANDOM}};
  r_501_0 = _RAND_3562[0:0];
  _RAND_3563 = {1{`RANDOM}};
  r_501_1 = _RAND_3563[0:0];
  _RAND_3564 = {1{`RANDOM}};
  r_502_0 = _RAND_3564[0:0];
  _RAND_3565 = {1{`RANDOM}};
  r_502_1 = _RAND_3565[0:0];
  _RAND_3566 = {1{`RANDOM}};
  r_503_0 = _RAND_3566[0:0];
  _RAND_3567 = {1{`RANDOM}};
  r_503_1 = _RAND_3567[0:0];
  _RAND_3568 = {1{`RANDOM}};
  r_504_0 = _RAND_3568[0:0];
  _RAND_3569 = {1{`RANDOM}};
  r_504_1 = _RAND_3569[0:0];
  _RAND_3570 = {1{`RANDOM}};
  r_505_0 = _RAND_3570[0:0];
  _RAND_3571 = {1{`RANDOM}};
  r_505_1 = _RAND_3571[0:0];
  _RAND_3572 = {1{`RANDOM}};
  r_506_0 = _RAND_3572[0:0];
  _RAND_3573 = {1{`RANDOM}};
  r_506_1 = _RAND_3573[0:0];
  _RAND_3574 = {1{`RANDOM}};
  r_507_0 = _RAND_3574[0:0];
  _RAND_3575 = {1{`RANDOM}};
  r_507_1 = _RAND_3575[0:0];
  _RAND_3576 = {1{`RANDOM}};
  r_508_0 = _RAND_3576[0:0];
  _RAND_3577 = {1{`RANDOM}};
  r_508_1 = _RAND_3577[0:0];
  _RAND_3578 = {1{`RANDOM}};
  r_509_0 = _RAND_3578[0:0];
  _RAND_3579 = {1{`RANDOM}};
  r_509_1 = _RAND_3579[0:0];
  _RAND_3580 = {1{`RANDOM}};
  r_510_0 = _RAND_3580[0:0];
  _RAND_3581 = {1{`RANDOM}};
  r_510_1 = _RAND_3581[0:0];
  _RAND_3582 = {1{`RANDOM}};
  r_511_0 = _RAND_3582[0:0];
  _RAND_3583 = {1{`RANDOM}};
  r_511_1 = _RAND_3583[0:0];
  _RAND_3584 = {1{`RANDOM}};
  r_512_0 = _RAND_3584[1:0];
  _RAND_3585 = {1{`RANDOM}};
  r_512_1 = _RAND_3585[1:0];
  _RAND_3586 = {1{`RANDOM}};
  r_513_0 = _RAND_3586[1:0];
  _RAND_3587 = {1{`RANDOM}};
  r_513_1 = _RAND_3587[1:0];
  _RAND_3588 = {1{`RANDOM}};
  r_514_0 = _RAND_3588[1:0];
  _RAND_3589 = {1{`RANDOM}};
  r_514_1 = _RAND_3589[1:0];
  _RAND_3590 = {1{`RANDOM}};
  r_515_0 = _RAND_3590[1:0];
  _RAND_3591 = {1{`RANDOM}};
  r_515_1 = _RAND_3591[1:0];
  _RAND_3592 = {1{`RANDOM}};
  r_516_0 = _RAND_3592[1:0];
  _RAND_3593 = {1{`RANDOM}};
  r_516_1 = _RAND_3593[1:0];
  _RAND_3594 = {1{`RANDOM}};
  r_517_0 = _RAND_3594[1:0];
  _RAND_3595 = {1{`RANDOM}};
  r_517_1 = _RAND_3595[1:0];
  _RAND_3596 = {1{`RANDOM}};
  r_518_0 = _RAND_3596[1:0];
  _RAND_3597 = {1{`RANDOM}};
  r_518_1 = _RAND_3597[1:0];
  _RAND_3598 = {1{`RANDOM}};
  r_519_0 = _RAND_3598[1:0];
  _RAND_3599 = {1{`RANDOM}};
  r_519_1 = _RAND_3599[1:0];
  _RAND_3600 = {1{`RANDOM}};
  r_520_0 = _RAND_3600[1:0];
  _RAND_3601 = {1{`RANDOM}};
  r_520_1 = _RAND_3601[1:0];
  _RAND_3602 = {1{`RANDOM}};
  r_521_0 = _RAND_3602[1:0];
  _RAND_3603 = {1{`RANDOM}};
  r_521_1 = _RAND_3603[1:0];
  _RAND_3604 = {1{`RANDOM}};
  r_522_0 = _RAND_3604[1:0];
  _RAND_3605 = {1{`RANDOM}};
  r_522_1 = _RAND_3605[1:0];
  _RAND_3606 = {1{`RANDOM}};
  r_523_0 = _RAND_3606[1:0];
  _RAND_3607 = {1{`RANDOM}};
  r_523_1 = _RAND_3607[1:0];
  _RAND_3608 = {1{`RANDOM}};
  r_524_0 = _RAND_3608[1:0];
  _RAND_3609 = {1{`RANDOM}};
  r_524_1 = _RAND_3609[1:0];
  _RAND_3610 = {1{`RANDOM}};
  r_525_0 = _RAND_3610[1:0];
  _RAND_3611 = {1{`RANDOM}};
  r_525_1 = _RAND_3611[1:0];
  _RAND_3612 = {1{`RANDOM}};
  r_526_0 = _RAND_3612[1:0];
  _RAND_3613 = {1{`RANDOM}};
  r_526_1 = _RAND_3613[1:0];
  _RAND_3614 = {1{`RANDOM}};
  r_527_0 = _RAND_3614[1:0];
  _RAND_3615 = {1{`RANDOM}};
  r_527_1 = _RAND_3615[1:0];
  _RAND_3616 = {1{`RANDOM}};
  r_528_0 = _RAND_3616[1:0];
  _RAND_3617 = {1{`RANDOM}};
  r_528_1 = _RAND_3617[1:0];
  _RAND_3618 = {1{`RANDOM}};
  r_529_0 = _RAND_3618[1:0];
  _RAND_3619 = {1{`RANDOM}};
  r_529_1 = _RAND_3619[1:0];
  _RAND_3620 = {1{`RANDOM}};
  r_530_0 = _RAND_3620[1:0];
  _RAND_3621 = {1{`RANDOM}};
  r_530_1 = _RAND_3621[1:0];
  _RAND_3622 = {1{`RANDOM}};
  r_531_0 = _RAND_3622[1:0];
  _RAND_3623 = {1{`RANDOM}};
  r_531_1 = _RAND_3623[1:0];
  _RAND_3624 = {1{`RANDOM}};
  r_532_0 = _RAND_3624[1:0];
  _RAND_3625 = {1{`RANDOM}};
  r_532_1 = _RAND_3625[1:0];
  _RAND_3626 = {1{`RANDOM}};
  r_533_0 = _RAND_3626[1:0];
  _RAND_3627 = {1{`RANDOM}};
  r_533_1 = _RAND_3627[1:0];
  _RAND_3628 = {1{`RANDOM}};
  r_534_0 = _RAND_3628[1:0];
  _RAND_3629 = {1{`RANDOM}};
  r_534_1 = _RAND_3629[1:0];
  _RAND_3630 = {1{`RANDOM}};
  r_535_0 = _RAND_3630[1:0];
  _RAND_3631 = {1{`RANDOM}};
  r_535_1 = _RAND_3631[1:0];
  _RAND_3632 = {1{`RANDOM}};
  r_536_0 = _RAND_3632[1:0];
  _RAND_3633 = {1{`RANDOM}};
  r_536_1 = _RAND_3633[1:0];
  _RAND_3634 = {1{`RANDOM}};
  r_537_0 = _RAND_3634[1:0];
  _RAND_3635 = {1{`RANDOM}};
  r_537_1 = _RAND_3635[1:0];
  _RAND_3636 = {1{`RANDOM}};
  r_538_0 = _RAND_3636[1:0];
  _RAND_3637 = {1{`RANDOM}};
  r_538_1 = _RAND_3637[1:0];
  _RAND_3638 = {1{`RANDOM}};
  r_539_0 = _RAND_3638[1:0];
  _RAND_3639 = {1{`RANDOM}};
  r_539_1 = _RAND_3639[1:0];
  _RAND_3640 = {1{`RANDOM}};
  r_540_0 = _RAND_3640[1:0];
  _RAND_3641 = {1{`RANDOM}};
  r_540_1 = _RAND_3641[1:0];
  _RAND_3642 = {1{`RANDOM}};
  r_541_0 = _RAND_3642[1:0];
  _RAND_3643 = {1{`RANDOM}};
  r_541_1 = _RAND_3643[1:0];
  _RAND_3644 = {1{`RANDOM}};
  r_542_0 = _RAND_3644[1:0];
  _RAND_3645 = {1{`RANDOM}};
  r_542_1 = _RAND_3645[1:0];
  _RAND_3646 = {1{`RANDOM}};
  r_543_0 = _RAND_3646[1:0];
  _RAND_3647 = {1{`RANDOM}};
  r_543_1 = _RAND_3647[1:0];
  _RAND_3648 = {1{`RANDOM}};
  r_544_0 = _RAND_3648[1:0];
  _RAND_3649 = {1{`RANDOM}};
  r_544_1 = _RAND_3649[1:0];
  _RAND_3650 = {1{`RANDOM}};
  r_545_0 = _RAND_3650[1:0];
  _RAND_3651 = {1{`RANDOM}};
  r_545_1 = _RAND_3651[1:0];
  _RAND_3652 = {1{`RANDOM}};
  r_546_0 = _RAND_3652[1:0];
  _RAND_3653 = {1{`RANDOM}};
  r_546_1 = _RAND_3653[1:0];
  _RAND_3654 = {1{`RANDOM}};
  r_547_0 = _RAND_3654[1:0];
  _RAND_3655 = {1{`RANDOM}};
  r_547_1 = _RAND_3655[1:0];
  _RAND_3656 = {1{`RANDOM}};
  r_548_0 = _RAND_3656[1:0];
  _RAND_3657 = {1{`RANDOM}};
  r_548_1 = _RAND_3657[1:0];
  _RAND_3658 = {1{`RANDOM}};
  r_549_0 = _RAND_3658[1:0];
  _RAND_3659 = {1{`RANDOM}};
  r_549_1 = _RAND_3659[1:0];
  _RAND_3660 = {1{`RANDOM}};
  r_550_0 = _RAND_3660[1:0];
  _RAND_3661 = {1{`RANDOM}};
  r_550_1 = _RAND_3661[1:0];
  _RAND_3662 = {1{`RANDOM}};
  r_551_0 = _RAND_3662[1:0];
  _RAND_3663 = {1{`RANDOM}};
  r_551_1 = _RAND_3663[1:0];
  _RAND_3664 = {1{`RANDOM}};
  r_552_0 = _RAND_3664[1:0];
  _RAND_3665 = {1{`RANDOM}};
  r_552_1 = _RAND_3665[1:0];
  _RAND_3666 = {1{`RANDOM}};
  r_553_0 = _RAND_3666[1:0];
  _RAND_3667 = {1{`RANDOM}};
  r_553_1 = _RAND_3667[1:0];
  _RAND_3668 = {1{`RANDOM}};
  r_554_0 = _RAND_3668[1:0];
  _RAND_3669 = {1{`RANDOM}};
  r_554_1 = _RAND_3669[1:0];
  _RAND_3670 = {1{`RANDOM}};
  r_555_0 = _RAND_3670[1:0];
  _RAND_3671 = {1{`RANDOM}};
  r_555_1 = _RAND_3671[1:0];
  _RAND_3672 = {1{`RANDOM}};
  r_556_0 = _RAND_3672[1:0];
  _RAND_3673 = {1{`RANDOM}};
  r_556_1 = _RAND_3673[1:0];
  _RAND_3674 = {1{`RANDOM}};
  r_557_0 = _RAND_3674[1:0];
  _RAND_3675 = {1{`RANDOM}};
  r_557_1 = _RAND_3675[1:0];
  _RAND_3676 = {1{`RANDOM}};
  r_558_0 = _RAND_3676[1:0];
  _RAND_3677 = {1{`RANDOM}};
  r_558_1 = _RAND_3677[1:0];
  _RAND_3678 = {1{`RANDOM}};
  r_559_0 = _RAND_3678[1:0];
  _RAND_3679 = {1{`RANDOM}};
  r_559_1 = _RAND_3679[1:0];
  _RAND_3680 = {1{`RANDOM}};
  r_560_0 = _RAND_3680[1:0];
  _RAND_3681 = {1{`RANDOM}};
  r_560_1 = _RAND_3681[1:0];
  _RAND_3682 = {1{`RANDOM}};
  r_561_0 = _RAND_3682[1:0];
  _RAND_3683 = {1{`RANDOM}};
  r_561_1 = _RAND_3683[1:0];
  _RAND_3684 = {1{`RANDOM}};
  r_562_0 = _RAND_3684[1:0];
  _RAND_3685 = {1{`RANDOM}};
  r_562_1 = _RAND_3685[1:0];
  _RAND_3686 = {1{`RANDOM}};
  r_563_0 = _RAND_3686[1:0];
  _RAND_3687 = {1{`RANDOM}};
  r_563_1 = _RAND_3687[1:0];
  _RAND_3688 = {1{`RANDOM}};
  r_564_0 = _RAND_3688[1:0];
  _RAND_3689 = {1{`RANDOM}};
  r_564_1 = _RAND_3689[1:0];
  _RAND_3690 = {1{`RANDOM}};
  r_565_0 = _RAND_3690[1:0];
  _RAND_3691 = {1{`RANDOM}};
  r_565_1 = _RAND_3691[1:0];
  _RAND_3692 = {1{`RANDOM}};
  r_566_0 = _RAND_3692[1:0];
  _RAND_3693 = {1{`RANDOM}};
  r_566_1 = _RAND_3693[1:0];
  _RAND_3694 = {1{`RANDOM}};
  r_567_0 = _RAND_3694[1:0];
  _RAND_3695 = {1{`RANDOM}};
  r_567_1 = _RAND_3695[1:0];
  _RAND_3696 = {1{`RANDOM}};
  r_568_0 = _RAND_3696[1:0];
  _RAND_3697 = {1{`RANDOM}};
  r_568_1 = _RAND_3697[1:0];
  _RAND_3698 = {1{`RANDOM}};
  r_569_0 = _RAND_3698[1:0];
  _RAND_3699 = {1{`RANDOM}};
  r_569_1 = _RAND_3699[1:0];
  _RAND_3700 = {1{`RANDOM}};
  r_570_0 = _RAND_3700[1:0];
  _RAND_3701 = {1{`RANDOM}};
  r_570_1 = _RAND_3701[1:0];
  _RAND_3702 = {1{`RANDOM}};
  r_571_0 = _RAND_3702[1:0];
  _RAND_3703 = {1{`RANDOM}};
  r_571_1 = _RAND_3703[1:0];
  _RAND_3704 = {1{`RANDOM}};
  r_572_0 = _RAND_3704[1:0];
  _RAND_3705 = {1{`RANDOM}};
  r_572_1 = _RAND_3705[1:0];
  _RAND_3706 = {1{`RANDOM}};
  r_573_0 = _RAND_3706[1:0];
  _RAND_3707 = {1{`RANDOM}};
  r_573_1 = _RAND_3707[1:0];
  _RAND_3708 = {1{`RANDOM}};
  r_574_0 = _RAND_3708[1:0];
  _RAND_3709 = {1{`RANDOM}};
  r_574_1 = _RAND_3709[1:0];
  _RAND_3710 = {1{`RANDOM}};
  r_575_0 = _RAND_3710[1:0];
  _RAND_3711 = {1{`RANDOM}};
  r_575_1 = _RAND_3711[1:0];
  _RAND_3712 = {1{`RANDOM}};
  r_576_0 = _RAND_3712[1:0];
  _RAND_3713 = {1{`RANDOM}};
  r_576_1 = _RAND_3713[1:0];
  _RAND_3714 = {1{`RANDOM}};
  r_577_0 = _RAND_3714[1:0];
  _RAND_3715 = {1{`RANDOM}};
  r_577_1 = _RAND_3715[1:0];
  _RAND_3716 = {1{`RANDOM}};
  r_578_0 = _RAND_3716[1:0];
  _RAND_3717 = {1{`RANDOM}};
  r_578_1 = _RAND_3717[1:0];
  _RAND_3718 = {1{`RANDOM}};
  r_579_0 = _RAND_3718[1:0];
  _RAND_3719 = {1{`RANDOM}};
  r_579_1 = _RAND_3719[1:0];
  _RAND_3720 = {1{`RANDOM}};
  r_580_0 = _RAND_3720[1:0];
  _RAND_3721 = {1{`RANDOM}};
  r_580_1 = _RAND_3721[1:0];
  _RAND_3722 = {1{`RANDOM}};
  r_581_0 = _RAND_3722[1:0];
  _RAND_3723 = {1{`RANDOM}};
  r_581_1 = _RAND_3723[1:0];
  _RAND_3724 = {1{`RANDOM}};
  r_582_0 = _RAND_3724[1:0];
  _RAND_3725 = {1{`RANDOM}};
  r_582_1 = _RAND_3725[1:0];
  _RAND_3726 = {1{`RANDOM}};
  r_583_0 = _RAND_3726[1:0];
  _RAND_3727 = {1{`RANDOM}};
  r_583_1 = _RAND_3727[1:0];
  _RAND_3728 = {1{`RANDOM}};
  r_584_0 = _RAND_3728[1:0];
  _RAND_3729 = {1{`RANDOM}};
  r_584_1 = _RAND_3729[1:0];
  _RAND_3730 = {1{`RANDOM}};
  r_585_0 = _RAND_3730[1:0];
  _RAND_3731 = {1{`RANDOM}};
  r_585_1 = _RAND_3731[1:0];
  _RAND_3732 = {1{`RANDOM}};
  r_586_0 = _RAND_3732[1:0];
  _RAND_3733 = {1{`RANDOM}};
  r_586_1 = _RAND_3733[1:0];
  _RAND_3734 = {1{`RANDOM}};
  r_587_0 = _RAND_3734[1:0];
  _RAND_3735 = {1{`RANDOM}};
  r_587_1 = _RAND_3735[1:0];
  _RAND_3736 = {1{`RANDOM}};
  r_588_0 = _RAND_3736[1:0];
  _RAND_3737 = {1{`RANDOM}};
  r_588_1 = _RAND_3737[1:0];
  _RAND_3738 = {1{`RANDOM}};
  r_589_0 = _RAND_3738[1:0];
  _RAND_3739 = {1{`RANDOM}};
  r_589_1 = _RAND_3739[1:0];
  _RAND_3740 = {1{`RANDOM}};
  r_590_0 = _RAND_3740[1:0];
  _RAND_3741 = {1{`RANDOM}};
  r_590_1 = _RAND_3741[1:0];
  _RAND_3742 = {1{`RANDOM}};
  r_591_0 = _RAND_3742[1:0];
  _RAND_3743 = {1{`RANDOM}};
  r_591_1 = _RAND_3743[1:0];
  _RAND_3744 = {1{`RANDOM}};
  r_592_0 = _RAND_3744[1:0];
  _RAND_3745 = {1{`RANDOM}};
  r_592_1 = _RAND_3745[1:0];
  _RAND_3746 = {1{`RANDOM}};
  r_593_0 = _RAND_3746[1:0];
  _RAND_3747 = {1{`RANDOM}};
  r_593_1 = _RAND_3747[1:0];
  _RAND_3748 = {1{`RANDOM}};
  r_594_0 = _RAND_3748[1:0];
  _RAND_3749 = {1{`RANDOM}};
  r_594_1 = _RAND_3749[1:0];
  _RAND_3750 = {1{`RANDOM}};
  r_595_0 = _RAND_3750[1:0];
  _RAND_3751 = {1{`RANDOM}};
  r_595_1 = _RAND_3751[1:0];
  _RAND_3752 = {1{`RANDOM}};
  r_596_0 = _RAND_3752[1:0];
  _RAND_3753 = {1{`RANDOM}};
  r_596_1 = _RAND_3753[1:0];
  _RAND_3754 = {1{`RANDOM}};
  r_597_0 = _RAND_3754[1:0];
  _RAND_3755 = {1{`RANDOM}};
  r_597_1 = _RAND_3755[1:0];
  _RAND_3756 = {1{`RANDOM}};
  r_598_0 = _RAND_3756[1:0];
  _RAND_3757 = {1{`RANDOM}};
  r_598_1 = _RAND_3757[1:0];
  _RAND_3758 = {1{`RANDOM}};
  r_599_0 = _RAND_3758[1:0];
  _RAND_3759 = {1{`RANDOM}};
  r_599_1 = _RAND_3759[1:0];
  _RAND_3760 = {1{`RANDOM}};
  r_600_0 = _RAND_3760[1:0];
  _RAND_3761 = {1{`RANDOM}};
  r_600_1 = _RAND_3761[1:0];
  _RAND_3762 = {1{`RANDOM}};
  r_601_0 = _RAND_3762[1:0];
  _RAND_3763 = {1{`RANDOM}};
  r_601_1 = _RAND_3763[1:0];
  _RAND_3764 = {1{`RANDOM}};
  r_602_0 = _RAND_3764[1:0];
  _RAND_3765 = {1{`RANDOM}};
  r_602_1 = _RAND_3765[1:0];
  _RAND_3766 = {1{`RANDOM}};
  r_603_0 = _RAND_3766[1:0];
  _RAND_3767 = {1{`RANDOM}};
  r_603_1 = _RAND_3767[1:0];
  _RAND_3768 = {1{`RANDOM}};
  r_604_0 = _RAND_3768[1:0];
  _RAND_3769 = {1{`RANDOM}};
  r_604_1 = _RAND_3769[1:0];
  _RAND_3770 = {1{`RANDOM}};
  r_605_0 = _RAND_3770[1:0];
  _RAND_3771 = {1{`RANDOM}};
  r_605_1 = _RAND_3771[1:0];
  _RAND_3772 = {1{`RANDOM}};
  r_606_0 = _RAND_3772[1:0];
  _RAND_3773 = {1{`RANDOM}};
  r_606_1 = _RAND_3773[1:0];
  _RAND_3774 = {1{`RANDOM}};
  r_607_0 = _RAND_3774[1:0];
  _RAND_3775 = {1{`RANDOM}};
  r_607_1 = _RAND_3775[1:0];
  _RAND_3776 = {1{`RANDOM}};
  r_608_0 = _RAND_3776[1:0];
  _RAND_3777 = {1{`RANDOM}};
  r_608_1 = _RAND_3777[1:0];
  _RAND_3778 = {1{`RANDOM}};
  r_609_0 = _RAND_3778[1:0];
  _RAND_3779 = {1{`RANDOM}};
  r_609_1 = _RAND_3779[1:0];
  _RAND_3780 = {1{`RANDOM}};
  r_610_0 = _RAND_3780[1:0];
  _RAND_3781 = {1{`RANDOM}};
  r_610_1 = _RAND_3781[1:0];
  _RAND_3782 = {1{`RANDOM}};
  r_611_0 = _RAND_3782[1:0];
  _RAND_3783 = {1{`RANDOM}};
  r_611_1 = _RAND_3783[1:0];
  _RAND_3784 = {1{`RANDOM}};
  r_612_0 = _RAND_3784[1:0];
  _RAND_3785 = {1{`RANDOM}};
  r_612_1 = _RAND_3785[1:0];
  _RAND_3786 = {1{`RANDOM}};
  r_613_0 = _RAND_3786[1:0];
  _RAND_3787 = {1{`RANDOM}};
  r_613_1 = _RAND_3787[1:0];
  _RAND_3788 = {1{`RANDOM}};
  r_614_0 = _RAND_3788[1:0];
  _RAND_3789 = {1{`RANDOM}};
  r_614_1 = _RAND_3789[1:0];
  _RAND_3790 = {1{`RANDOM}};
  r_615_0 = _RAND_3790[1:0];
  _RAND_3791 = {1{`RANDOM}};
  r_615_1 = _RAND_3791[1:0];
  _RAND_3792 = {1{`RANDOM}};
  r_616_0 = _RAND_3792[1:0];
  _RAND_3793 = {1{`RANDOM}};
  r_616_1 = _RAND_3793[1:0];
  _RAND_3794 = {1{`RANDOM}};
  r_617_0 = _RAND_3794[1:0];
  _RAND_3795 = {1{`RANDOM}};
  r_617_1 = _RAND_3795[1:0];
  _RAND_3796 = {1{`RANDOM}};
  r_618_0 = _RAND_3796[1:0];
  _RAND_3797 = {1{`RANDOM}};
  r_618_1 = _RAND_3797[1:0];
  _RAND_3798 = {1{`RANDOM}};
  r_619_0 = _RAND_3798[1:0];
  _RAND_3799 = {1{`RANDOM}};
  r_619_1 = _RAND_3799[1:0];
  _RAND_3800 = {1{`RANDOM}};
  r_620_0 = _RAND_3800[1:0];
  _RAND_3801 = {1{`RANDOM}};
  r_620_1 = _RAND_3801[1:0];
  _RAND_3802 = {1{`RANDOM}};
  r_621_0 = _RAND_3802[1:0];
  _RAND_3803 = {1{`RANDOM}};
  r_621_1 = _RAND_3803[1:0];
  _RAND_3804 = {1{`RANDOM}};
  r_622_0 = _RAND_3804[1:0];
  _RAND_3805 = {1{`RANDOM}};
  r_622_1 = _RAND_3805[1:0];
  _RAND_3806 = {1{`RANDOM}};
  r_623_0 = _RAND_3806[1:0];
  _RAND_3807 = {1{`RANDOM}};
  r_623_1 = _RAND_3807[1:0];
  _RAND_3808 = {1{`RANDOM}};
  r_624_0 = _RAND_3808[1:0];
  _RAND_3809 = {1{`RANDOM}};
  r_624_1 = _RAND_3809[1:0];
  _RAND_3810 = {1{`RANDOM}};
  r_625_0 = _RAND_3810[1:0];
  _RAND_3811 = {1{`RANDOM}};
  r_625_1 = _RAND_3811[1:0];
  _RAND_3812 = {1{`RANDOM}};
  r_626_0 = _RAND_3812[1:0];
  _RAND_3813 = {1{`RANDOM}};
  r_626_1 = _RAND_3813[1:0];
  _RAND_3814 = {1{`RANDOM}};
  r_627_0 = _RAND_3814[1:0];
  _RAND_3815 = {1{`RANDOM}};
  r_627_1 = _RAND_3815[1:0];
  _RAND_3816 = {1{`RANDOM}};
  r_628_0 = _RAND_3816[1:0];
  _RAND_3817 = {1{`RANDOM}};
  r_628_1 = _RAND_3817[1:0];
  _RAND_3818 = {1{`RANDOM}};
  r_629_0 = _RAND_3818[1:0];
  _RAND_3819 = {1{`RANDOM}};
  r_629_1 = _RAND_3819[1:0];
  _RAND_3820 = {1{`RANDOM}};
  r_630_0 = _RAND_3820[1:0];
  _RAND_3821 = {1{`RANDOM}};
  r_630_1 = _RAND_3821[1:0];
  _RAND_3822 = {1{`RANDOM}};
  r_631_0 = _RAND_3822[1:0];
  _RAND_3823 = {1{`RANDOM}};
  r_631_1 = _RAND_3823[1:0];
  _RAND_3824 = {1{`RANDOM}};
  r_632_0 = _RAND_3824[1:0];
  _RAND_3825 = {1{`RANDOM}};
  r_632_1 = _RAND_3825[1:0];
  _RAND_3826 = {1{`RANDOM}};
  r_633_0 = _RAND_3826[1:0];
  _RAND_3827 = {1{`RANDOM}};
  r_633_1 = _RAND_3827[1:0];
  _RAND_3828 = {1{`RANDOM}};
  r_634_0 = _RAND_3828[1:0];
  _RAND_3829 = {1{`RANDOM}};
  r_634_1 = _RAND_3829[1:0];
  _RAND_3830 = {1{`RANDOM}};
  r_635_0 = _RAND_3830[1:0];
  _RAND_3831 = {1{`RANDOM}};
  r_635_1 = _RAND_3831[1:0];
  _RAND_3832 = {1{`RANDOM}};
  r_636_0 = _RAND_3832[1:0];
  _RAND_3833 = {1{`RANDOM}};
  r_636_1 = _RAND_3833[1:0];
  _RAND_3834 = {1{`RANDOM}};
  r_637_0 = _RAND_3834[1:0];
  _RAND_3835 = {1{`RANDOM}};
  r_637_1 = _RAND_3835[1:0];
  _RAND_3836 = {1{`RANDOM}};
  r_638_0 = _RAND_3836[1:0];
  _RAND_3837 = {1{`RANDOM}};
  r_638_1 = _RAND_3837[1:0];
  _RAND_3838 = {1{`RANDOM}};
  r_639_0 = _RAND_3838[1:0];
  _RAND_3839 = {1{`RANDOM}};
  r_639_1 = _RAND_3839[1:0];
  _RAND_3840 = {1{`RANDOM}};
  r_640_0 = _RAND_3840[1:0];
  _RAND_3841 = {1{`RANDOM}};
  r_640_1 = _RAND_3841[1:0];
  _RAND_3842 = {1{`RANDOM}};
  r_641_0 = _RAND_3842[1:0];
  _RAND_3843 = {1{`RANDOM}};
  r_641_1 = _RAND_3843[1:0];
  _RAND_3844 = {1{`RANDOM}};
  r_642_0 = _RAND_3844[1:0];
  _RAND_3845 = {1{`RANDOM}};
  r_642_1 = _RAND_3845[1:0];
  _RAND_3846 = {1{`RANDOM}};
  r_643_0 = _RAND_3846[1:0];
  _RAND_3847 = {1{`RANDOM}};
  r_643_1 = _RAND_3847[1:0];
  _RAND_3848 = {1{`RANDOM}};
  r_644_0 = _RAND_3848[1:0];
  _RAND_3849 = {1{`RANDOM}};
  r_644_1 = _RAND_3849[1:0];
  _RAND_3850 = {1{`RANDOM}};
  r_645_0 = _RAND_3850[1:0];
  _RAND_3851 = {1{`RANDOM}};
  r_645_1 = _RAND_3851[1:0];
  _RAND_3852 = {1{`RANDOM}};
  r_646_0 = _RAND_3852[1:0];
  _RAND_3853 = {1{`RANDOM}};
  r_646_1 = _RAND_3853[1:0];
  _RAND_3854 = {1{`RANDOM}};
  r_647_0 = _RAND_3854[1:0];
  _RAND_3855 = {1{`RANDOM}};
  r_647_1 = _RAND_3855[1:0];
  _RAND_3856 = {1{`RANDOM}};
  r_648_0 = _RAND_3856[1:0];
  _RAND_3857 = {1{`RANDOM}};
  r_648_1 = _RAND_3857[1:0];
  _RAND_3858 = {1{`RANDOM}};
  r_649_0 = _RAND_3858[1:0];
  _RAND_3859 = {1{`RANDOM}};
  r_649_1 = _RAND_3859[1:0];
  _RAND_3860 = {1{`RANDOM}};
  r_650_0 = _RAND_3860[1:0];
  _RAND_3861 = {1{`RANDOM}};
  r_650_1 = _RAND_3861[1:0];
  _RAND_3862 = {1{`RANDOM}};
  r_651_0 = _RAND_3862[1:0];
  _RAND_3863 = {1{`RANDOM}};
  r_651_1 = _RAND_3863[1:0];
  _RAND_3864 = {1{`RANDOM}};
  r_652_0 = _RAND_3864[1:0];
  _RAND_3865 = {1{`RANDOM}};
  r_652_1 = _RAND_3865[1:0];
  _RAND_3866 = {1{`RANDOM}};
  r_653_0 = _RAND_3866[1:0];
  _RAND_3867 = {1{`RANDOM}};
  r_653_1 = _RAND_3867[1:0];
  _RAND_3868 = {1{`RANDOM}};
  r_654_0 = _RAND_3868[1:0];
  _RAND_3869 = {1{`RANDOM}};
  r_654_1 = _RAND_3869[1:0];
  _RAND_3870 = {1{`RANDOM}};
  r_655_0 = _RAND_3870[1:0];
  _RAND_3871 = {1{`RANDOM}};
  r_655_1 = _RAND_3871[1:0];
  _RAND_3872 = {1{`RANDOM}};
  r_656_0 = _RAND_3872[1:0];
  _RAND_3873 = {1{`RANDOM}};
  r_656_1 = _RAND_3873[1:0];
  _RAND_3874 = {1{`RANDOM}};
  r_657_0 = _RAND_3874[1:0];
  _RAND_3875 = {1{`RANDOM}};
  r_657_1 = _RAND_3875[1:0];
  _RAND_3876 = {1{`RANDOM}};
  r_658_0 = _RAND_3876[1:0];
  _RAND_3877 = {1{`RANDOM}};
  r_658_1 = _RAND_3877[1:0];
  _RAND_3878 = {1{`RANDOM}};
  r_659_0 = _RAND_3878[1:0];
  _RAND_3879 = {1{`RANDOM}};
  r_659_1 = _RAND_3879[1:0];
  _RAND_3880 = {1{`RANDOM}};
  r_660_0 = _RAND_3880[1:0];
  _RAND_3881 = {1{`RANDOM}};
  r_660_1 = _RAND_3881[1:0];
  _RAND_3882 = {1{`RANDOM}};
  r_661_0 = _RAND_3882[1:0];
  _RAND_3883 = {1{`RANDOM}};
  r_661_1 = _RAND_3883[1:0];
  _RAND_3884 = {1{`RANDOM}};
  r_662_0 = _RAND_3884[1:0];
  _RAND_3885 = {1{`RANDOM}};
  r_662_1 = _RAND_3885[1:0];
  _RAND_3886 = {1{`RANDOM}};
  r_663_0 = _RAND_3886[1:0];
  _RAND_3887 = {1{`RANDOM}};
  r_663_1 = _RAND_3887[1:0];
  _RAND_3888 = {1{`RANDOM}};
  r_664_0 = _RAND_3888[1:0];
  _RAND_3889 = {1{`RANDOM}};
  r_664_1 = _RAND_3889[1:0];
  _RAND_3890 = {1{`RANDOM}};
  r_665_0 = _RAND_3890[1:0];
  _RAND_3891 = {1{`RANDOM}};
  r_665_1 = _RAND_3891[1:0];
  _RAND_3892 = {1{`RANDOM}};
  r_666_0 = _RAND_3892[1:0];
  _RAND_3893 = {1{`RANDOM}};
  r_666_1 = _RAND_3893[1:0];
  _RAND_3894 = {1{`RANDOM}};
  r_667_0 = _RAND_3894[1:0];
  _RAND_3895 = {1{`RANDOM}};
  r_667_1 = _RAND_3895[1:0];
  _RAND_3896 = {1{`RANDOM}};
  r_668_0 = _RAND_3896[1:0];
  _RAND_3897 = {1{`RANDOM}};
  r_668_1 = _RAND_3897[1:0];
  _RAND_3898 = {1{`RANDOM}};
  r_669_0 = _RAND_3898[1:0];
  _RAND_3899 = {1{`RANDOM}};
  r_669_1 = _RAND_3899[1:0];
  _RAND_3900 = {1{`RANDOM}};
  r_670_0 = _RAND_3900[1:0];
  _RAND_3901 = {1{`RANDOM}};
  r_670_1 = _RAND_3901[1:0];
  _RAND_3902 = {1{`RANDOM}};
  r_671_0 = _RAND_3902[1:0];
  _RAND_3903 = {1{`RANDOM}};
  r_671_1 = _RAND_3903[1:0];
  _RAND_3904 = {1{`RANDOM}};
  r_672_0 = _RAND_3904[1:0];
  _RAND_3905 = {1{`RANDOM}};
  r_672_1 = _RAND_3905[1:0];
  _RAND_3906 = {1{`RANDOM}};
  r_673_0 = _RAND_3906[1:0];
  _RAND_3907 = {1{`RANDOM}};
  r_673_1 = _RAND_3907[1:0];
  _RAND_3908 = {1{`RANDOM}};
  r_674_0 = _RAND_3908[1:0];
  _RAND_3909 = {1{`RANDOM}};
  r_674_1 = _RAND_3909[1:0];
  _RAND_3910 = {1{`RANDOM}};
  r_675_0 = _RAND_3910[1:0];
  _RAND_3911 = {1{`RANDOM}};
  r_675_1 = _RAND_3911[1:0];
  _RAND_3912 = {1{`RANDOM}};
  r_676_0 = _RAND_3912[1:0];
  _RAND_3913 = {1{`RANDOM}};
  r_676_1 = _RAND_3913[1:0];
  _RAND_3914 = {1{`RANDOM}};
  r_677_0 = _RAND_3914[1:0];
  _RAND_3915 = {1{`RANDOM}};
  r_677_1 = _RAND_3915[1:0];
  _RAND_3916 = {1{`RANDOM}};
  r_678_0 = _RAND_3916[1:0];
  _RAND_3917 = {1{`RANDOM}};
  r_678_1 = _RAND_3917[1:0];
  _RAND_3918 = {1{`RANDOM}};
  r_679_0 = _RAND_3918[1:0];
  _RAND_3919 = {1{`RANDOM}};
  r_679_1 = _RAND_3919[1:0];
  _RAND_3920 = {1{`RANDOM}};
  r_680_0 = _RAND_3920[1:0];
  _RAND_3921 = {1{`RANDOM}};
  r_680_1 = _RAND_3921[1:0];
  _RAND_3922 = {1{`RANDOM}};
  r_681_0 = _RAND_3922[1:0];
  _RAND_3923 = {1{`RANDOM}};
  r_681_1 = _RAND_3923[1:0];
  _RAND_3924 = {1{`RANDOM}};
  r_682_0 = _RAND_3924[1:0];
  _RAND_3925 = {1{`RANDOM}};
  r_682_1 = _RAND_3925[1:0];
  _RAND_3926 = {1{`RANDOM}};
  r_683_0 = _RAND_3926[1:0];
  _RAND_3927 = {1{`RANDOM}};
  r_683_1 = _RAND_3927[1:0];
  _RAND_3928 = {1{`RANDOM}};
  r_684_0 = _RAND_3928[1:0];
  _RAND_3929 = {1{`RANDOM}};
  r_684_1 = _RAND_3929[1:0];
  _RAND_3930 = {1{`RANDOM}};
  r_685_0 = _RAND_3930[1:0];
  _RAND_3931 = {1{`RANDOM}};
  r_685_1 = _RAND_3931[1:0];
  _RAND_3932 = {1{`RANDOM}};
  r_686_0 = _RAND_3932[1:0];
  _RAND_3933 = {1{`RANDOM}};
  r_686_1 = _RAND_3933[1:0];
  _RAND_3934 = {1{`RANDOM}};
  r_687_0 = _RAND_3934[1:0];
  _RAND_3935 = {1{`RANDOM}};
  r_687_1 = _RAND_3935[1:0];
  _RAND_3936 = {1{`RANDOM}};
  r_688_0 = _RAND_3936[1:0];
  _RAND_3937 = {1{`RANDOM}};
  r_688_1 = _RAND_3937[1:0];
  _RAND_3938 = {1{`RANDOM}};
  r_689_0 = _RAND_3938[1:0];
  _RAND_3939 = {1{`RANDOM}};
  r_689_1 = _RAND_3939[1:0];
  _RAND_3940 = {1{`RANDOM}};
  r_690_0 = _RAND_3940[1:0];
  _RAND_3941 = {1{`RANDOM}};
  r_690_1 = _RAND_3941[1:0];
  _RAND_3942 = {1{`RANDOM}};
  r_691_0 = _RAND_3942[1:0];
  _RAND_3943 = {1{`RANDOM}};
  r_691_1 = _RAND_3943[1:0];
  _RAND_3944 = {1{`RANDOM}};
  r_692_0 = _RAND_3944[1:0];
  _RAND_3945 = {1{`RANDOM}};
  r_692_1 = _RAND_3945[1:0];
  _RAND_3946 = {1{`RANDOM}};
  r_693_0 = _RAND_3946[1:0];
  _RAND_3947 = {1{`RANDOM}};
  r_693_1 = _RAND_3947[1:0];
  _RAND_3948 = {1{`RANDOM}};
  r_694_0 = _RAND_3948[1:0];
  _RAND_3949 = {1{`RANDOM}};
  r_694_1 = _RAND_3949[1:0];
  _RAND_3950 = {1{`RANDOM}};
  r_695_0 = _RAND_3950[1:0];
  _RAND_3951 = {1{`RANDOM}};
  r_695_1 = _RAND_3951[1:0];
  _RAND_3952 = {1{`RANDOM}};
  r_696_0 = _RAND_3952[1:0];
  _RAND_3953 = {1{`RANDOM}};
  r_696_1 = _RAND_3953[1:0];
  _RAND_3954 = {1{`RANDOM}};
  r_697_0 = _RAND_3954[1:0];
  _RAND_3955 = {1{`RANDOM}};
  r_697_1 = _RAND_3955[1:0];
  _RAND_3956 = {1{`RANDOM}};
  r_698_0 = _RAND_3956[1:0];
  _RAND_3957 = {1{`RANDOM}};
  r_698_1 = _RAND_3957[1:0];
  _RAND_3958 = {1{`RANDOM}};
  r_699_0 = _RAND_3958[1:0];
  _RAND_3959 = {1{`RANDOM}};
  r_699_1 = _RAND_3959[1:0];
  _RAND_3960 = {1{`RANDOM}};
  r_700_0 = _RAND_3960[1:0];
  _RAND_3961 = {1{`RANDOM}};
  r_700_1 = _RAND_3961[1:0];
  _RAND_3962 = {1{`RANDOM}};
  r_701_0 = _RAND_3962[1:0];
  _RAND_3963 = {1{`RANDOM}};
  r_701_1 = _RAND_3963[1:0];
  _RAND_3964 = {1{`RANDOM}};
  r_702_0 = _RAND_3964[1:0];
  _RAND_3965 = {1{`RANDOM}};
  r_702_1 = _RAND_3965[1:0];
  _RAND_3966 = {1{`RANDOM}};
  r_703_0 = _RAND_3966[1:0];
  _RAND_3967 = {1{`RANDOM}};
  r_703_1 = _RAND_3967[1:0];
  _RAND_3968 = {1{`RANDOM}};
  r_704_0 = _RAND_3968[1:0];
  _RAND_3969 = {1{`RANDOM}};
  r_704_1 = _RAND_3969[1:0];
  _RAND_3970 = {1{`RANDOM}};
  r_705_0 = _RAND_3970[1:0];
  _RAND_3971 = {1{`RANDOM}};
  r_705_1 = _RAND_3971[1:0];
  _RAND_3972 = {1{`RANDOM}};
  r_706_0 = _RAND_3972[1:0];
  _RAND_3973 = {1{`RANDOM}};
  r_706_1 = _RAND_3973[1:0];
  _RAND_3974 = {1{`RANDOM}};
  r_707_0 = _RAND_3974[1:0];
  _RAND_3975 = {1{`RANDOM}};
  r_707_1 = _RAND_3975[1:0];
  _RAND_3976 = {1{`RANDOM}};
  r_708_0 = _RAND_3976[1:0];
  _RAND_3977 = {1{`RANDOM}};
  r_708_1 = _RAND_3977[1:0];
  _RAND_3978 = {1{`RANDOM}};
  r_709_0 = _RAND_3978[1:0];
  _RAND_3979 = {1{`RANDOM}};
  r_709_1 = _RAND_3979[1:0];
  _RAND_3980 = {1{`RANDOM}};
  r_710_0 = _RAND_3980[1:0];
  _RAND_3981 = {1{`RANDOM}};
  r_710_1 = _RAND_3981[1:0];
  _RAND_3982 = {1{`RANDOM}};
  r_711_0 = _RAND_3982[1:0];
  _RAND_3983 = {1{`RANDOM}};
  r_711_1 = _RAND_3983[1:0];
  _RAND_3984 = {1{`RANDOM}};
  r_712_0 = _RAND_3984[1:0];
  _RAND_3985 = {1{`RANDOM}};
  r_712_1 = _RAND_3985[1:0];
  _RAND_3986 = {1{`RANDOM}};
  r_713_0 = _RAND_3986[1:0];
  _RAND_3987 = {1{`RANDOM}};
  r_713_1 = _RAND_3987[1:0];
  _RAND_3988 = {1{`RANDOM}};
  r_714_0 = _RAND_3988[1:0];
  _RAND_3989 = {1{`RANDOM}};
  r_714_1 = _RAND_3989[1:0];
  _RAND_3990 = {1{`RANDOM}};
  r_715_0 = _RAND_3990[1:0];
  _RAND_3991 = {1{`RANDOM}};
  r_715_1 = _RAND_3991[1:0];
  _RAND_3992 = {1{`RANDOM}};
  r_716_0 = _RAND_3992[1:0];
  _RAND_3993 = {1{`RANDOM}};
  r_716_1 = _RAND_3993[1:0];
  _RAND_3994 = {1{`RANDOM}};
  r_717_0 = _RAND_3994[1:0];
  _RAND_3995 = {1{`RANDOM}};
  r_717_1 = _RAND_3995[1:0];
  _RAND_3996 = {1{`RANDOM}};
  r_718_0 = _RAND_3996[1:0];
  _RAND_3997 = {1{`RANDOM}};
  r_718_1 = _RAND_3997[1:0];
  _RAND_3998 = {1{`RANDOM}};
  r_719_0 = _RAND_3998[1:0];
  _RAND_3999 = {1{`RANDOM}};
  r_719_1 = _RAND_3999[1:0];
  _RAND_4000 = {1{`RANDOM}};
  r_720_0 = _RAND_4000[1:0];
  _RAND_4001 = {1{`RANDOM}};
  r_720_1 = _RAND_4001[1:0];
  _RAND_4002 = {1{`RANDOM}};
  r_721_0 = _RAND_4002[1:0];
  _RAND_4003 = {1{`RANDOM}};
  r_721_1 = _RAND_4003[1:0];
  _RAND_4004 = {1{`RANDOM}};
  r_722_0 = _RAND_4004[1:0];
  _RAND_4005 = {1{`RANDOM}};
  r_722_1 = _RAND_4005[1:0];
  _RAND_4006 = {1{`RANDOM}};
  r_723_0 = _RAND_4006[1:0];
  _RAND_4007 = {1{`RANDOM}};
  r_723_1 = _RAND_4007[1:0];
  _RAND_4008 = {1{`RANDOM}};
  r_724_0 = _RAND_4008[1:0];
  _RAND_4009 = {1{`RANDOM}};
  r_724_1 = _RAND_4009[1:0];
  _RAND_4010 = {1{`RANDOM}};
  r_725_0 = _RAND_4010[1:0];
  _RAND_4011 = {1{`RANDOM}};
  r_725_1 = _RAND_4011[1:0];
  _RAND_4012 = {1{`RANDOM}};
  r_726_0 = _RAND_4012[1:0];
  _RAND_4013 = {1{`RANDOM}};
  r_726_1 = _RAND_4013[1:0];
  _RAND_4014 = {1{`RANDOM}};
  r_727_0 = _RAND_4014[1:0];
  _RAND_4015 = {1{`RANDOM}};
  r_727_1 = _RAND_4015[1:0];
  _RAND_4016 = {1{`RANDOM}};
  r_728_0 = _RAND_4016[1:0];
  _RAND_4017 = {1{`RANDOM}};
  r_728_1 = _RAND_4017[1:0];
  _RAND_4018 = {1{`RANDOM}};
  r_729_0 = _RAND_4018[1:0];
  _RAND_4019 = {1{`RANDOM}};
  r_729_1 = _RAND_4019[1:0];
  _RAND_4020 = {1{`RANDOM}};
  r_730_0 = _RAND_4020[1:0];
  _RAND_4021 = {1{`RANDOM}};
  r_730_1 = _RAND_4021[1:0];
  _RAND_4022 = {1{`RANDOM}};
  r_731_0 = _RAND_4022[1:0];
  _RAND_4023 = {1{`RANDOM}};
  r_731_1 = _RAND_4023[1:0];
  _RAND_4024 = {1{`RANDOM}};
  r_732_0 = _RAND_4024[1:0];
  _RAND_4025 = {1{`RANDOM}};
  r_732_1 = _RAND_4025[1:0];
  _RAND_4026 = {1{`RANDOM}};
  r_733_0 = _RAND_4026[1:0];
  _RAND_4027 = {1{`RANDOM}};
  r_733_1 = _RAND_4027[1:0];
  _RAND_4028 = {1{`RANDOM}};
  r_734_0 = _RAND_4028[1:0];
  _RAND_4029 = {1{`RANDOM}};
  r_734_1 = _RAND_4029[1:0];
  _RAND_4030 = {1{`RANDOM}};
  r_735_0 = _RAND_4030[1:0];
  _RAND_4031 = {1{`RANDOM}};
  r_735_1 = _RAND_4031[1:0];
  _RAND_4032 = {1{`RANDOM}};
  r_736_0 = _RAND_4032[1:0];
  _RAND_4033 = {1{`RANDOM}};
  r_736_1 = _RAND_4033[1:0];
  _RAND_4034 = {1{`RANDOM}};
  r_737_0 = _RAND_4034[1:0];
  _RAND_4035 = {1{`RANDOM}};
  r_737_1 = _RAND_4035[1:0];
  _RAND_4036 = {1{`RANDOM}};
  r_738_0 = _RAND_4036[1:0];
  _RAND_4037 = {1{`RANDOM}};
  r_738_1 = _RAND_4037[1:0];
  _RAND_4038 = {1{`RANDOM}};
  r_739_0 = _RAND_4038[1:0];
  _RAND_4039 = {1{`RANDOM}};
  r_739_1 = _RAND_4039[1:0];
  _RAND_4040 = {1{`RANDOM}};
  r_740_0 = _RAND_4040[1:0];
  _RAND_4041 = {1{`RANDOM}};
  r_740_1 = _RAND_4041[1:0];
  _RAND_4042 = {1{`RANDOM}};
  r_741_0 = _RAND_4042[1:0];
  _RAND_4043 = {1{`RANDOM}};
  r_741_1 = _RAND_4043[1:0];
  _RAND_4044 = {1{`RANDOM}};
  r_742_0 = _RAND_4044[1:0];
  _RAND_4045 = {1{`RANDOM}};
  r_742_1 = _RAND_4045[1:0];
  _RAND_4046 = {1{`RANDOM}};
  r_743_0 = _RAND_4046[1:0];
  _RAND_4047 = {1{`RANDOM}};
  r_743_1 = _RAND_4047[1:0];
  _RAND_4048 = {1{`RANDOM}};
  r_744_0 = _RAND_4048[1:0];
  _RAND_4049 = {1{`RANDOM}};
  r_744_1 = _RAND_4049[1:0];
  _RAND_4050 = {1{`RANDOM}};
  r_745_0 = _RAND_4050[1:0];
  _RAND_4051 = {1{`RANDOM}};
  r_745_1 = _RAND_4051[1:0];
  _RAND_4052 = {1{`RANDOM}};
  r_746_0 = _RAND_4052[1:0];
  _RAND_4053 = {1{`RANDOM}};
  r_746_1 = _RAND_4053[1:0];
  _RAND_4054 = {1{`RANDOM}};
  r_747_0 = _RAND_4054[1:0];
  _RAND_4055 = {1{`RANDOM}};
  r_747_1 = _RAND_4055[1:0];
  _RAND_4056 = {1{`RANDOM}};
  r_748_0 = _RAND_4056[1:0];
  _RAND_4057 = {1{`RANDOM}};
  r_748_1 = _RAND_4057[1:0];
  _RAND_4058 = {1{`RANDOM}};
  r_749_0 = _RAND_4058[1:0];
  _RAND_4059 = {1{`RANDOM}};
  r_749_1 = _RAND_4059[1:0];
  _RAND_4060 = {1{`RANDOM}};
  r_750_0 = _RAND_4060[1:0];
  _RAND_4061 = {1{`RANDOM}};
  r_750_1 = _RAND_4061[1:0];
  _RAND_4062 = {1{`RANDOM}};
  r_751_0 = _RAND_4062[1:0];
  _RAND_4063 = {1{`RANDOM}};
  r_751_1 = _RAND_4063[1:0];
  _RAND_4064 = {1{`RANDOM}};
  r_752_0 = _RAND_4064[1:0];
  _RAND_4065 = {1{`RANDOM}};
  r_752_1 = _RAND_4065[1:0];
  _RAND_4066 = {1{`RANDOM}};
  r_753_0 = _RAND_4066[1:0];
  _RAND_4067 = {1{`RANDOM}};
  r_753_1 = _RAND_4067[1:0];
  _RAND_4068 = {1{`RANDOM}};
  r_754_0 = _RAND_4068[1:0];
  _RAND_4069 = {1{`RANDOM}};
  r_754_1 = _RAND_4069[1:0];
  _RAND_4070 = {1{`RANDOM}};
  r_755_0 = _RAND_4070[1:0];
  _RAND_4071 = {1{`RANDOM}};
  r_755_1 = _RAND_4071[1:0];
  _RAND_4072 = {1{`RANDOM}};
  r_756_0 = _RAND_4072[1:0];
  _RAND_4073 = {1{`RANDOM}};
  r_756_1 = _RAND_4073[1:0];
  _RAND_4074 = {1{`RANDOM}};
  r_757_0 = _RAND_4074[1:0];
  _RAND_4075 = {1{`RANDOM}};
  r_757_1 = _RAND_4075[1:0];
  _RAND_4076 = {1{`RANDOM}};
  r_758_0 = _RAND_4076[1:0];
  _RAND_4077 = {1{`RANDOM}};
  r_758_1 = _RAND_4077[1:0];
  _RAND_4078 = {1{`RANDOM}};
  r_759_0 = _RAND_4078[1:0];
  _RAND_4079 = {1{`RANDOM}};
  r_759_1 = _RAND_4079[1:0];
  _RAND_4080 = {1{`RANDOM}};
  r_760_0 = _RAND_4080[1:0];
  _RAND_4081 = {1{`RANDOM}};
  r_760_1 = _RAND_4081[1:0];
  _RAND_4082 = {1{`RANDOM}};
  r_761_0 = _RAND_4082[1:0];
  _RAND_4083 = {1{`RANDOM}};
  r_761_1 = _RAND_4083[1:0];
  _RAND_4084 = {1{`RANDOM}};
  r_762_0 = _RAND_4084[1:0];
  _RAND_4085 = {1{`RANDOM}};
  r_762_1 = _RAND_4085[1:0];
  _RAND_4086 = {1{`RANDOM}};
  r_763_0 = _RAND_4086[1:0];
  _RAND_4087 = {1{`RANDOM}};
  r_763_1 = _RAND_4087[1:0];
  _RAND_4088 = {1{`RANDOM}};
  r_764_0 = _RAND_4088[1:0];
  _RAND_4089 = {1{`RANDOM}};
  r_764_1 = _RAND_4089[1:0];
  _RAND_4090 = {1{`RANDOM}};
  r_765_0 = _RAND_4090[1:0];
  _RAND_4091 = {1{`RANDOM}};
  r_765_1 = _RAND_4091[1:0];
  _RAND_4092 = {1{`RANDOM}};
  r_766_0 = _RAND_4092[1:0];
  _RAND_4093 = {1{`RANDOM}};
  r_766_1 = _RAND_4093[1:0];
  _RAND_4094 = {1{`RANDOM}};
  r_767_0 = _RAND_4094[1:0];
  _RAND_4095 = {1{`RANDOM}};
  r_767_1 = _RAND_4095[1:0];
  _RAND_4096 = {1{`RANDOM}};
  r_768_0 = _RAND_4096[0:0];
  _RAND_4097 = {1{`RANDOM}};
  r_768_1 = _RAND_4097[0:0];
  _RAND_4098 = {1{`RANDOM}};
  r_769_0 = _RAND_4098[0:0];
  _RAND_4099 = {1{`RANDOM}};
  r_769_1 = _RAND_4099[0:0];
  _RAND_4100 = {1{`RANDOM}};
  r_770_0 = _RAND_4100[0:0];
  _RAND_4101 = {1{`RANDOM}};
  r_770_1 = _RAND_4101[0:0];
  _RAND_4102 = {1{`RANDOM}};
  r_771_0 = _RAND_4102[0:0];
  _RAND_4103 = {1{`RANDOM}};
  r_771_1 = _RAND_4103[0:0];
  _RAND_4104 = {1{`RANDOM}};
  r_772_0 = _RAND_4104[0:0];
  _RAND_4105 = {1{`RANDOM}};
  r_772_1 = _RAND_4105[0:0];
  _RAND_4106 = {1{`RANDOM}};
  r_773_0 = _RAND_4106[0:0];
  _RAND_4107 = {1{`RANDOM}};
  r_773_1 = _RAND_4107[0:0];
  _RAND_4108 = {1{`RANDOM}};
  r_774_0 = _RAND_4108[0:0];
  _RAND_4109 = {1{`RANDOM}};
  r_774_1 = _RAND_4109[0:0];
  _RAND_4110 = {1{`RANDOM}};
  r_775_0 = _RAND_4110[0:0];
  _RAND_4111 = {1{`RANDOM}};
  r_775_1 = _RAND_4111[0:0];
  _RAND_4112 = {1{`RANDOM}};
  r_776_0 = _RAND_4112[0:0];
  _RAND_4113 = {1{`RANDOM}};
  r_776_1 = _RAND_4113[0:0];
  _RAND_4114 = {1{`RANDOM}};
  r_777_0 = _RAND_4114[0:0];
  _RAND_4115 = {1{`RANDOM}};
  r_777_1 = _RAND_4115[0:0];
  _RAND_4116 = {1{`RANDOM}};
  r_778_0 = _RAND_4116[0:0];
  _RAND_4117 = {1{`RANDOM}};
  r_778_1 = _RAND_4117[0:0];
  _RAND_4118 = {1{`RANDOM}};
  r_779_0 = _RAND_4118[0:0];
  _RAND_4119 = {1{`RANDOM}};
  r_779_1 = _RAND_4119[0:0];
  _RAND_4120 = {1{`RANDOM}};
  r_780_0 = _RAND_4120[0:0];
  _RAND_4121 = {1{`RANDOM}};
  r_780_1 = _RAND_4121[0:0];
  _RAND_4122 = {1{`RANDOM}};
  r_781_0 = _RAND_4122[0:0];
  _RAND_4123 = {1{`RANDOM}};
  r_781_1 = _RAND_4123[0:0];
  _RAND_4124 = {1{`RANDOM}};
  r_782_0 = _RAND_4124[0:0];
  _RAND_4125 = {1{`RANDOM}};
  r_782_1 = _RAND_4125[0:0];
  _RAND_4126 = {1{`RANDOM}};
  r_783_0 = _RAND_4126[0:0];
  _RAND_4127 = {1{`RANDOM}};
  r_783_1 = _RAND_4127[0:0];
  _RAND_4128 = {1{`RANDOM}};
  r_784_0 = _RAND_4128[0:0];
  _RAND_4129 = {1{`RANDOM}};
  r_784_1 = _RAND_4129[0:0];
  _RAND_4130 = {1{`RANDOM}};
  r_785_0 = _RAND_4130[0:0];
  _RAND_4131 = {1{`RANDOM}};
  r_785_1 = _RAND_4131[0:0];
  _RAND_4132 = {1{`RANDOM}};
  r_786_0 = _RAND_4132[0:0];
  _RAND_4133 = {1{`RANDOM}};
  r_786_1 = _RAND_4133[0:0];
  _RAND_4134 = {1{`RANDOM}};
  r_787_0 = _RAND_4134[0:0];
  _RAND_4135 = {1{`RANDOM}};
  r_787_1 = _RAND_4135[0:0];
  _RAND_4136 = {1{`RANDOM}};
  r_788_0 = _RAND_4136[0:0];
  _RAND_4137 = {1{`RANDOM}};
  r_788_1 = _RAND_4137[0:0];
  _RAND_4138 = {1{`RANDOM}};
  r_789_0 = _RAND_4138[0:0];
  _RAND_4139 = {1{`RANDOM}};
  r_789_1 = _RAND_4139[0:0];
  _RAND_4140 = {1{`RANDOM}};
  r_790_0 = _RAND_4140[0:0];
  _RAND_4141 = {1{`RANDOM}};
  r_790_1 = _RAND_4141[0:0];
  _RAND_4142 = {1{`RANDOM}};
  r_791_0 = _RAND_4142[0:0];
  _RAND_4143 = {1{`RANDOM}};
  r_791_1 = _RAND_4143[0:0];
  _RAND_4144 = {1{`RANDOM}};
  r_792_0 = _RAND_4144[0:0];
  _RAND_4145 = {1{`RANDOM}};
  r_792_1 = _RAND_4145[0:0];
  _RAND_4146 = {1{`RANDOM}};
  r_793_0 = _RAND_4146[0:0];
  _RAND_4147 = {1{`RANDOM}};
  r_793_1 = _RAND_4147[0:0];
  _RAND_4148 = {1{`RANDOM}};
  r_794_0 = _RAND_4148[0:0];
  _RAND_4149 = {1{`RANDOM}};
  r_794_1 = _RAND_4149[0:0];
  _RAND_4150 = {1{`RANDOM}};
  r_795_0 = _RAND_4150[0:0];
  _RAND_4151 = {1{`RANDOM}};
  r_795_1 = _RAND_4151[0:0];
  _RAND_4152 = {1{`RANDOM}};
  r_796_0 = _RAND_4152[0:0];
  _RAND_4153 = {1{`RANDOM}};
  r_796_1 = _RAND_4153[0:0];
  _RAND_4154 = {1{`RANDOM}};
  r_797_0 = _RAND_4154[0:0];
  _RAND_4155 = {1{`RANDOM}};
  r_797_1 = _RAND_4155[0:0];
  _RAND_4156 = {1{`RANDOM}};
  r_798_0 = _RAND_4156[0:0];
  _RAND_4157 = {1{`RANDOM}};
  r_798_1 = _RAND_4157[0:0];
  _RAND_4158 = {1{`RANDOM}};
  r_799_0 = _RAND_4158[0:0];
  _RAND_4159 = {1{`RANDOM}};
  r_799_1 = _RAND_4159[0:0];
  _RAND_4160 = {1{`RANDOM}};
  r_800_0 = _RAND_4160[0:0];
  _RAND_4161 = {1{`RANDOM}};
  r_800_1 = _RAND_4161[0:0];
  _RAND_4162 = {1{`RANDOM}};
  r_801_0 = _RAND_4162[0:0];
  _RAND_4163 = {1{`RANDOM}};
  r_801_1 = _RAND_4163[0:0];
  _RAND_4164 = {1{`RANDOM}};
  r_802_0 = _RAND_4164[0:0];
  _RAND_4165 = {1{`RANDOM}};
  r_802_1 = _RAND_4165[0:0];
  _RAND_4166 = {1{`RANDOM}};
  r_803_0 = _RAND_4166[0:0];
  _RAND_4167 = {1{`RANDOM}};
  r_803_1 = _RAND_4167[0:0];
  _RAND_4168 = {1{`RANDOM}};
  r_804_0 = _RAND_4168[0:0];
  _RAND_4169 = {1{`RANDOM}};
  r_804_1 = _RAND_4169[0:0];
  _RAND_4170 = {1{`RANDOM}};
  r_805_0 = _RAND_4170[0:0];
  _RAND_4171 = {1{`RANDOM}};
  r_805_1 = _RAND_4171[0:0];
  _RAND_4172 = {1{`RANDOM}};
  r_806_0 = _RAND_4172[0:0];
  _RAND_4173 = {1{`RANDOM}};
  r_806_1 = _RAND_4173[0:0];
  _RAND_4174 = {1{`RANDOM}};
  r_807_0 = _RAND_4174[0:0];
  _RAND_4175 = {1{`RANDOM}};
  r_807_1 = _RAND_4175[0:0];
  _RAND_4176 = {1{`RANDOM}};
  r_808_0 = _RAND_4176[0:0];
  _RAND_4177 = {1{`RANDOM}};
  r_808_1 = _RAND_4177[0:0];
  _RAND_4178 = {1{`RANDOM}};
  r_809_0 = _RAND_4178[0:0];
  _RAND_4179 = {1{`RANDOM}};
  r_809_1 = _RAND_4179[0:0];
  _RAND_4180 = {1{`RANDOM}};
  r_810_0 = _RAND_4180[0:0];
  _RAND_4181 = {1{`RANDOM}};
  r_810_1 = _RAND_4181[0:0];
  _RAND_4182 = {1{`RANDOM}};
  r_811_0 = _RAND_4182[0:0];
  _RAND_4183 = {1{`RANDOM}};
  r_811_1 = _RAND_4183[0:0];
  _RAND_4184 = {1{`RANDOM}};
  r_812_0 = _RAND_4184[0:0];
  _RAND_4185 = {1{`RANDOM}};
  r_812_1 = _RAND_4185[0:0];
  _RAND_4186 = {1{`RANDOM}};
  r_813_0 = _RAND_4186[0:0];
  _RAND_4187 = {1{`RANDOM}};
  r_813_1 = _RAND_4187[0:0];
  _RAND_4188 = {1{`RANDOM}};
  r_814_0 = _RAND_4188[0:0];
  _RAND_4189 = {1{`RANDOM}};
  r_814_1 = _RAND_4189[0:0];
  _RAND_4190 = {1{`RANDOM}};
  r_815_0 = _RAND_4190[0:0];
  _RAND_4191 = {1{`RANDOM}};
  r_815_1 = _RAND_4191[0:0];
  _RAND_4192 = {1{`RANDOM}};
  r_816_0 = _RAND_4192[0:0];
  _RAND_4193 = {1{`RANDOM}};
  r_816_1 = _RAND_4193[0:0];
  _RAND_4194 = {1{`RANDOM}};
  r_817_0 = _RAND_4194[0:0];
  _RAND_4195 = {1{`RANDOM}};
  r_817_1 = _RAND_4195[0:0];
  _RAND_4196 = {1{`RANDOM}};
  r_818_0 = _RAND_4196[0:0];
  _RAND_4197 = {1{`RANDOM}};
  r_818_1 = _RAND_4197[0:0];
  _RAND_4198 = {1{`RANDOM}};
  r_819_0 = _RAND_4198[0:0];
  _RAND_4199 = {1{`RANDOM}};
  r_819_1 = _RAND_4199[0:0];
  _RAND_4200 = {1{`RANDOM}};
  r_820_0 = _RAND_4200[0:0];
  _RAND_4201 = {1{`RANDOM}};
  r_820_1 = _RAND_4201[0:0];
  _RAND_4202 = {1{`RANDOM}};
  r_821_0 = _RAND_4202[0:0];
  _RAND_4203 = {1{`RANDOM}};
  r_821_1 = _RAND_4203[0:0];
  _RAND_4204 = {1{`RANDOM}};
  r_822_0 = _RAND_4204[0:0];
  _RAND_4205 = {1{`RANDOM}};
  r_822_1 = _RAND_4205[0:0];
  _RAND_4206 = {1{`RANDOM}};
  r_823_0 = _RAND_4206[0:0];
  _RAND_4207 = {1{`RANDOM}};
  r_823_1 = _RAND_4207[0:0];
  _RAND_4208 = {1{`RANDOM}};
  r_824_0 = _RAND_4208[0:0];
  _RAND_4209 = {1{`RANDOM}};
  r_824_1 = _RAND_4209[0:0];
  _RAND_4210 = {1{`RANDOM}};
  r_825_0 = _RAND_4210[0:0];
  _RAND_4211 = {1{`RANDOM}};
  r_825_1 = _RAND_4211[0:0];
  _RAND_4212 = {1{`RANDOM}};
  r_826_0 = _RAND_4212[0:0];
  _RAND_4213 = {1{`RANDOM}};
  r_826_1 = _RAND_4213[0:0];
  _RAND_4214 = {1{`RANDOM}};
  r_827_0 = _RAND_4214[0:0];
  _RAND_4215 = {1{`RANDOM}};
  r_827_1 = _RAND_4215[0:0];
  _RAND_4216 = {1{`RANDOM}};
  r_828_0 = _RAND_4216[0:0];
  _RAND_4217 = {1{`RANDOM}};
  r_828_1 = _RAND_4217[0:0];
  _RAND_4218 = {1{`RANDOM}};
  r_829_0 = _RAND_4218[0:0];
  _RAND_4219 = {1{`RANDOM}};
  r_829_1 = _RAND_4219[0:0];
  _RAND_4220 = {1{`RANDOM}};
  r_830_0 = _RAND_4220[0:0];
  _RAND_4221 = {1{`RANDOM}};
  r_830_1 = _RAND_4221[0:0];
  _RAND_4222 = {1{`RANDOM}};
  r_831_0 = _RAND_4222[0:0];
  _RAND_4223 = {1{`RANDOM}};
  r_831_1 = _RAND_4223[0:0];
  _RAND_4224 = {1{`RANDOM}};
  r_832_0 = _RAND_4224[0:0];
  _RAND_4225 = {1{`RANDOM}};
  r_832_1 = _RAND_4225[0:0];
  _RAND_4226 = {1{`RANDOM}};
  r_833_0 = _RAND_4226[0:0];
  _RAND_4227 = {1{`RANDOM}};
  r_833_1 = _RAND_4227[0:0];
  _RAND_4228 = {1{`RANDOM}};
  r_834_0 = _RAND_4228[0:0];
  _RAND_4229 = {1{`RANDOM}};
  r_834_1 = _RAND_4229[0:0];
  _RAND_4230 = {1{`RANDOM}};
  r_835_0 = _RAND_4230[0:0];
  _RAND_4231 = {1{`RANDOM}};
  r_835_1 = _RAND_4231[0:0];
  _RAND_4232 = {1{`RANDOM}};
  r_836_0 = _RAND_4232[0:0];
  _RAND_4233 = {1{`RANDOM}};
  r_836_1 = _RAND_4233[0:0];
  _RAND_4234 = {1{`RANDOM}};
  r_837_0 = _RAND_4234[0:0];
  _RAND_4235 = {1{`RANDOM}};
  r_837_1 = _RAND_4235[0:0];
  _RAND_4236 = {1{`RANDOM}};
  r_838_0 = _RAND_4236[0:0];
  _RAND_4237 = {1{`RANDOM}};
  r_838_1 = _RAND_4237[0:0];
  _RAND_4238 = {1{`RANDOM}};
  r_839_0 = _RAND_4238[0:0];
  _RAND_4239 = {1{`RANDOM}};
  r_839_1 = _RAND_4239[0:0];
  _RAND_4240 = {1{`RANDOM}};
  r_840_0 = _RAND_4240[0:0];
  _RAND_4241 = {1{`RANDOM}};
  r_840_1 = _RAND_4241[0:0];
  _RAND_4242 = {1{`RANDOM}};
  r_841_0 = _RAND_4242[0:0];
  _RAND_4243 = {1{`RANDOM}};
  r_841_1 = _RAND_4243[0:0];
  _RAND_4244 = {1{`RANDOM}};
  r_842_0 = _RAND_4244[0:0];
  _RAND_4245 = {1{`RANDOM}};
  r_842_1 = _RAND_4245[0:0];
  _RAND_4246 = {1{`RANDOM}};
  r_843_0 = _RAND_4246[0:0];
  _RAND_4247 = {1{`RANDOM}};
  r_843_1 = _RAND_4247[0:0];
  _RAND_4248 = {1{`RANDOM}};
  r_844_0 = _RAND_4248[0:0];
  _RAND_4249 = {1{`RANDOM}};
  r_844_1 = _RAND_4249[0:0];
  _RAND_4250 = {1{`RANDOM}};
  r_845_0 = _RAND_4250[0:0];
  _RAND_4251 = {1{`RANDOM}};
  r_845_1 = _RAND_4251[0:0];
  _RAND_4252 = {1{`RANDOM}};
  r_846_0 = _RAND_4252[0:0];
  _RAND_4253 = {1{`RANDOM}};
  r_846_1 = _RAND_4253[0:0];
  _RAND_4254 = {1{`RANDOM}};
  r_847_0 = _RAND_4254[0:0];
  _RAND_4255 = {1{`RANDOM}};
  r_847_1 = _RAND_4255[0:0];
  _RAND_4256 = {1{`RANDOM}};
  r_848_0 = _RAND_4256[0:0];
  _RAND_4257 = {1{`RANDOM}};
  r_848_1 = _RAND_4257[0:0];
  _RAND_4258 = {1{`RANDOM}};
  r_849_0 = _RAND_4258[0:0];
  _RAND_4259 = {1{`RANDOM}};
  r_849_1 = _RAND_4259[0:0];
  _RAND_4260 = {1{`RANDOM}};
  r_850_0 = _RAND_4260[0:0];
  _RAND_4261 = {1{`RANDOM}};
  r_850_1 = _RAND_4261[0:0];
  _RAND_4262 = {1{`RANDOM}};
  r_851_0 = _RAND_4262[0:0];
  _RAND_4263 = {1{`RANDOM}};
  r_851_1 = _RAND_4263[0:0];
  _RAND_4264 = {1{`RANDOM}};
  r_852_0 = _RAND_4264[0:0];
  _RAND_4265 = {1{`RANDOM}};
  r_852_1 = _RAND_4265[0:0];
  _RAND_4266 = {1{`RANDOM}};
  r_853_0 = _RAND_4266[0:0];
  _RAND_4267 = {1{`RANDOM}};
  r_853_1 = _RAND_4267[0:0];
  _RAND_4268 = {1{`RANDOM}};
  r_854_0 = _RAND_4268[0:0];
  _RAND_4269 = {1{`RANDOM}};
  r_854_1 = _RAND_4269[0:0];
  _RAND_4270 = {1{`RANDOM}};
  r_855_0 = _RAND_4270[0:0];
  _RAND_4271 = {1{`RANDOM}};
  r_855_1 = _RAND_4271[0:0];
  _RAND_4272 = {1{`RANDOM}};
  r_856_0 = _RAND_4272[0:0];
  _RAND_4273 = {1{`RANDOM}};
  r_856_1 = _RAND_4273[0:0];
  _RAND_4274 = {1{`RANDOM}};
  r_857_0 = _RAND_4274[0:0];
  _RAND_4275 = {1{`RANDOM}};
  r_857_1 = _RAND_4275[0:0];
  _RAND_4276 = {1{`RANDOM}};
  r_858_0 = _RAND_4276[0:0];
  _RAND_4277 = {1{`RANDOM}};
  r_858_1 = _RAND_4277[0:0];
  _RAND_4278 = {1{`RANDOM}};
  r_859_0 = _RAND_4278[0:0];
  _RAND_4279 = {1{`RANDOM}};
  r_859_1 = _RAND_4279[0:0];
  _RAND_4280 = {1{`RANDOM}};
  r_860_0 = _RAND_4280[0:0];
  _RAND_4281 = {1{`RANDOM}};
  r_860_1 = _RAND_4281[0:0];
  _RAND_4282 = {1{`RANDOM}};
  r_861_0 = _RAND_4282[0:0];
  _RAND_4283 = {1{`RANDOM}};
  r_861_1 = _RAND_4283[0:0];
  _RAND_4284 = {1{`RANDOM}};
  r_862_0 = _RAND_4284[0:0];
  _RAND_4285 = {1{`RANDOM}};
  r_862_1 = _RAND_4285[0:0];
  _RAND_4286 = {1{`RANDOM}};
  r_863_0 = _RAND_4286[0:0];
  _RAND_4287 = {1{`RANDOM}};
  r_863_1 = _RAND_4287[0:0];
  _RAND_4288 = {1{`RANDOM}};
  r_864_0 = _RAND_4288[0:0];
  _RAND_4289 = {1{`RANDOM}};
  r_864_1 = _RAND_4289[0:0];
  _RAND_4290 = {1{`RANDOM}};
  r_865_0 = _RAND_4290[0:0];
  _RAND_4291 = {1{`RANDOM}};
  r_865_1 = _RAND_4291[0:0];
  _RAND_4292 = {1{`RANDOM}};
  r_866_0 = _RAND_4292[0:0];
  _RAND_4293 = {1{`RANDOM}};
  r_866_1 = _RAND_4293[0:0];
  _RAND_4294 = {1{`RANDOM}};
  r_867_0 = _RAND_4294[0:0];
  _RAND_4295 = {1{`RANDOM}};
  r_867_1 = _RAND_4295[0:0];
  _RAND_4296 = {1{`RANDOM}};
  r_868_0 = _RAND_4296[0:0];
  _RAND_4297 = {1{`RANDOM}};
  r_868_1 = _RAND_4297[0:0];
  _RAND_4298 = {1{`RANDOM}};
  r_869_0 = _RAND_4298[0:0];
  _RAND_4299 = {1{`RANDOM}};
  r_869_1 = _RAND_4299[0:0];
  _RAND_4300 = {1{`RANDOM}};
  r_870_0 = _RAND_4300[0:0];
  _RAND_4301 = {1{`RANDOM}};
  r_870_1 = _RAND_4301[0:0];
  _RAND_4302 = {1{`RANDOM}};
  r_871_0 = _RAND_4302[0:0];
  _RAND_4303 = {1{`RANDOM}};
  r_871_1 = _RAND_4303[0:0];
  _RAND_4304 = {1{`RANDOM}};
  r_872_0 = _RAND_4304[0:0];
  _RAND_4305 = {1{`RANDOM}};
  r_872_1 = _RAND_4305[0:0];
  _RAND_4306 = {1{`RANDOM}};
  r_873_0 = _RAND_4306[0:0];
  _RAND_4307 = {1{`RANDOM}};
  r_873_1 = _RAND_4307[0:0];
  _RAND_4308 = {1{`RANDOM}};
  r_874_0 = _RAND_4308[0:0];
  _RAND_4309 = {1{`RANDOM}};
  r_874_1 = _RAND_4309[0:0];
  _RAND_4310 = {1{`RANDOM}};
  r_875_0 = _RAND_4310[0:0];
  _RAND_4311 = {1{`RANDOM}};
  r_875_1 = _RAND_4311[0:0];
  _RAND_4312 = {1{`RANDOM}};
  r_876_0 = _RAND_4312[0:0];
  _RAND_4313 = {1{`RANDOM}};
  r_876_1 = _RAND_4313[0:0];
  _RAND_4314 = {1{`RANDOM}};
  r_877_0 = _RAND_4314[0:0];
  _RAND_4315 = {1{`RANDOM}};
  r_877_1 = _RAND_4315[0:0];
  _RAND_4316 = {1{`RANDOM}};
  r_878_0 = _RAND_4316[0:0];
  _RAND_4317 = {1{`RANDOM}};
  r_878_1 = _RAND_4317[0:0];
  _RAND_4318 = {1{`RANDOM}};
  r_879_0 = _RAND_4318[0:0];
  _RAND_4319 = {1{`RANDOM}};
  r_879_1 = _RAND_4319[0:0];
  _RAND_4320 = {1{`RANDOM}};
  r_880_0 = _RAND_4320[0:0];
  _RAND_4321 = {1{`RANDOM}};
  r_880_1 = _RAND_4321[0:0];
  _RAND_4322 = {1{`RANDOM}};
  r_881_0 = _RAND_4322[0:0];
  _RAND_4323 = {1{`RANDOM}};
  r_881_1 = _RAND_4323[0:0];
  _RAND_4324 = {1{`RANDOM}};
  r_882_0 = _RAND_4324[0:0];
  _RAND_4325 = {1{`RANDOM}};
  r_882_1 = _RAND_4325[0:0];
  _RAND_4326 = {1{`RANDOM}};
  r_883_0 = _RAND_4326[0:0];
  _RAND_4327 = {1{`RANDOM}};
  r_883_1 = _RAND_4327[0:0];
  _RAND_4328 = {1{`RANDOM}};
  r_884_0 = _RAND_4328[0:0];
  _RAND_4329 = {1{`RANDOM}};
  r_884_1 = _RAND_4329[0:0];
  _RAND_4330 = {1{`RANDOM}};
  r_885_0 = _RAND_4330[0:0];
  _RAND_4331 = {1{`RANDOM}};
  r_885_1 = _RAND_4331[0:0];
  _RAND_4332 = {1{`RANDOM}};
  r_886_0 = _RAND_4332[0:0];
  _RAND_4333 = {1{`RANDOM}};
  r_886_1 = _RAND_4333[0:0];
  _RAND_4334 = {1{`RANDOM}};
  r_887_0 = _RAND_4334[0:0];
  _RAND_4335 = {1{`RANDOM}};
  r_887_1 = _RAND_4335[0:0];
  _RAND_4336 = {1{`RANDOM}};
  r_888_0 = _RAND_4336[0:0];
  _RAND_4337 = {1{`RANDOM}};
  r_888_1 = _RAND_4337[0:0];
  _RAND_4338 = {1{`RANDOM}};
  r_889_0 = _RAND_4338[0:0];
  _RAND_4339 = {1{`RANDOM}};
  r_889_1 = _RAND_4339[0:0];
  _RAND_4340 = {1{`RANDOM}};
  r_890_0 = _RAND_4340[0:0];
  _RAND_4341 = {1{`RANDOM}};
  r_890_1 = _RAND_4341[0:0];
  _RAND_4342 = {1{`RANDOM}};
  r_891_0 = _RAND_4342[0:0];
  _RAND_4343 = {1{`RANDOM}};
  r_891_1 = _RAND_4343[0:0];
  _RAND_4344 = {1{`RANDOM}};
  r_892_0 = _RAND_4344[0:0];
  _RAND_4345 = {1{`RANDOM}};
  r_892_1 = _RAND_4345[0:0];
  _RAND_4346 = {1{`RANDOM}};
  r_893_0 = _RAND_4346[0:0];
  _RAND_4347 = {1{`RANDOM}};
  r_893_1 = _RAND_4347[0:0];
  _RAND_4348 = {1{`RANDOM}};
  r_894_0 = _RAND_4348[0:0];
  _RAND_4349 = {1{`RANDOM}};
  r_894_1 = _RAND_4349[0:0];
  _RAND_4350 = {1{`RANDOM}};
  r_895_0 = _RAND_4350[0:0];
  _RAND_4351 = {1{`RANDOM}};
  r_895_1 = _RAND_4351[0:0];
  _RAND_4352 = {1{`RANDOM}};
  r_896_0 = _RAND_4352[0:0];
  _RAND_4353 = {1{`RANDOM}};
  r_896_1 = _RAND_4353[0:0];
  _RAND_4354 = {1{`RANDOM}};
  r_897_0 = _RAND_4354[0:0];
  _RAND_4355 = {1{`RANDOM}};
  r_897_1 = _RAND_4355[0:0];
  _RAND_4356 = {1{`RANDOM}};
  r_898_0 = _RAND_4356[0:0];
  _RAND_4357 = {1{`RANDOM}};
  r_898_1 = _RAND_4357[0:0];
  _RAND_4358 = {1{`RANDOM}};
  r_899_0 = _RAND_4358[0:0];
  _RAND_4359 = {1{`RANDOM}};
  r_899_1 = _RAND_4359[0:0];
  _RAND_4360 = {1{`RANDOM}};
  r_900_0 = _RAND_4360[0:0];
  _RAND_4361 = {1{`RANDOM}};
  r_900_1 = _RAND_4361[0:0];
  _RAND_4362 = {1{`RANDOM}};
  r_901_0 = _RAND_4362[0:0];
  _RAND_4363 = {1{`RANDOM}};
  r_901_1 = _RAND_4363[0:0];
  _RAND_4364 = {1{`RANDOM}};
  r_902_0 = _RAND_4364[0:0];
  _RAND_4365 = {1{`RANDOM}};
  r_902_1 = _RAND_4365[0:0];
  _RAND_4366 = {1{`RANDOM}};
  r_903_0 = _RAND_4366[0:0];
  _RAND_4367 = {1{`RANDOM}};
  r_903_1 = _RAND_4367[0:0];
  _RAND_4368 = {1{`RANDOM}};
  r_904_0 = _RAND_4368[0:0];
  _RAND_4369 = {1{`RANDOM}};
  r_904_1 = _RAND_4369[0:0];
  _RAND_4370 = {1{`RANDOM}};
  r_905_0 = _RAND_4370[0:0];
  _RAND_4371 = {1{`RANDOM}};
  r_905_1 = _RAND_4371[0:0];
  _RAND_4372 = {1{`RANDOM}};
  r_906_0 = _RAND_4372[0:0];
  _RAND_4373 = {1{`RANDOM}};
  r_906_1 = _RAND_4373[0:0];
  _RAND_4374 = {1{`RANDOM}};
  r_907_0 = _RAND_4374[0:0];
  _RAND_4375 = {1{`RANDOM}};
  r_907_1 = _RAND_4375[0:0];
  _RAND_4376 = {1{`RANDOM}};
  r_908_0 = _RAND_4376[0:0];
  _RAND_4377 = {1{`RANDOM}};
  r_908_1 = _RAND_4377[0:0];
  _RAND_4378 = {1{`RANDOM}};
  r_909_0 = _RAND_4378[0:0];
  _RAND_4379 = {1{`RANDOM}};
  r_909_1 = _RAND_4379[0:0];
  _RAND_4380 = {1{`RANDOM}};
  r_910_0 = _RAND_4380[0:0];
  _RAND_4381 = {1{`RANDOM}};
  r_910_1 = _RAND_4381[0:0];
  _RAND_4382 = {1{`RANDOM}};
  r_911_0 = _RAND_4382[0:0];
  _RAND_4383 = {1{`RANDOM}};
  r_911_1 = _RAND_4383[0:0];
  _RAND_4384 = {1{`RANDOM}};
  r_912_0 = _RAND_4384[0:0];
  _RAND_4385 = {1{`RANDOM}};
  r_912_1 = _RAND_4385[0:0];
  _RAND_4386 = {1{`RANDOM}};
  r_913_0 = _RAND_4386[0:0];
  _RAND_4387 = {1{`RANDOM}};
  r_913_1 = _RAND_4387[0:0];
  _RAND_4388 = {1{`RANDOM}};
  r_914_0 = _RAND_4388[0:0];
  _RAND_4389 = {1{`RANDOM}};
  r_914_1 = _RAND_4389[0:0];
  _RAND_4390 = {1{`RANDOM}};
  r_915_0 = _RAND_4390[0:0];
  _RAND_4391 = {1{`RANDOM}};
  r_915_1 = _RAND_4391[0:0];
  _RAND_4392 = {1{`RANDOM}};
  r_916_0 = _RAND_4392[0:0];
  _RAND_4393 = {1{`RANDOM}};
  r_916_1 = _RAND_4393[0:0];
  _RAND_4394 = {1{`RANDOM}};
  r_917_0 = _RAND_4394[0:0];
  _RAND_4395 = {1{`RANDOM}};
  r_917_1 = _RAND_4395[0:0];
  _RAND_4396 = {1{`RANDOM}};
  r_918_0 = _RAND_4396[0:0];
  _RAND_4397 = {1{`RANDOM}};
  r_918_1 = _RAND_4397[0:0];
  _RAND_4398 = {1{`RANDOM}};
  r_919_0 = _RAND_4398[0:0];
  _RAND_4399 = {1{`RANDOM}};
  r_919_1 = _RAND_4399[0:0];
  _RAND_4400 = {1{`RANDOM}};
  r_920_0 = _RAND_4400[0:0];
  _RAND_4401 = {1{`RANDOM}};
  r_920_1 = _RAND_4401[0:0];
  _RAND_4402 = {1{`RANDOM}};
  r_921_0 = _RAND_4402[0:0];
  _RAND_4403 = {1{`RANDOM}};
  r_921_1 = _RAND_4403[0:0];
  _RAND_4404 = {1{`RANDOM}};
  r_922_0 = _RAND_4404[0:0];
  _RAND_4405 = {1{`RANDOM}};
  r_922_1 = _RAND_4405[0:0];
  _RAND_4406 = {1{`RANDOM}};
  r_923_0 = _RAND_4406[0:0];
  _RAND_4407 = {1{`RANDOM}};
  r_923_1 = _RAND_4407[0:0];
  _RAND_4408 = {1{`RANDOM}};
  r_924_0 = _RAND_4408[0:0];
  _RAND_4409 = {1{`RANDOM}};
  r_924_1 = _RAND_4409[0:0];
  _RAND_4410 = {1{`RANDOM}};
  r_925_0 = _RAND_4410[0:0];
  _RAND_4411 = {1{`RANDOM}};
  r_925_1 = _RAND_4411[0:0];
  _RAND_4412 = {1{`RANDOM}};
  r_926_0 = _RAND_4412[0:0];
  _RAND_4413 = {1{`RANDOM}};
  r_926_1 = _RAND_4413[0:0];
  _RAND_4414 = {1{`RANDOM}};
  r_927_0 = _RAND_4414[0:0];
  _RAND_4415 = {1{`RANDOM}};
  r_927_1 = _RAND_4415[0:0];
  _RAND_4416 = {1{`RANDOM}};
  r_928_0 = _RAND_4416[0:0];
  _RAND_4417 = {1{`RANDOM}};
  r_928_1 = _RAND_4417[0:0];
  _RAND_4418 = {1{`RANDOM}};
  r_929_0 = _RAND_4418[0:0];
  _RAND_4419 = {1{`RANDOM}};
  r_929_1 = _RAND_4419[0:0];
  _RAND_4420 = {1{`RANDOM}};
  r_930_0 = _RAND_4420[0:0];
  _RAND_4421 = {1{`RANDOM}};
  r_930_1 = _RAND_4421[0:0];
  _RAND_4422 = {1{`RANDOM}};
  r_931_0 = _RAND_4422[0:0];
  _RAND_4423 = {1{`RANDOM}};
  r_931_1 = _RAND_4423[0:0];
  _RAND_4424 = {1{`RANDOM}};
  r_932_0 = _RAND_4424[0:0];
  _RAND_4425 = {1{`RANDOM}};
  r_932_1 = _RAND_4425[0:0];
  _RAND_4426 = {1{`RANDOM}};
  r_933_0 = _RAND_4426[0:0];
  _RAND_4427 = {1{`RANDOM}};
  r_933_1 = _RAND_4427[0:0];
  _RAND_4428 = {1{`RANDOM}};
  r_934_0 = _RAND_4428[0:0];
  _RAND_4429 = {1{`RANDOM}};
  r_934_1 = _RAND_4429[0:0];
  _RAND_4430 = {1{`RANDOM}};
  r_935_0 = _RAND_4430[0:0];
  _RAND_4431 = {1{`RANDOM}};
  r_935_1 = _RAND_4431[0:0];
  _RAND_4432 = {1{`RANDOM}};
  r_936_0 = _RAND_4432[0:0];
  _RAND_4433 = {1{`RANDOM}};
  r_936_1 = _RAND_4433[0:0];
  _RAND_4434 = {1{`RANDOM}};
  r_937_0 = _RAND_4434[0:0];
  _RAND_4435 = {1{`RANDOM}};
  r_937_1 = _RAND_4435[0:0];
  _RAND_4436 = {1{`RANDOM}};
  r_938_0 = _RAND_4436[0:0];
  _RAND_4437 = {1{`RANDOM}};
  r_938_1 = _RAND_4437[0:0];
  _RAND_4438 = {1{`RANDOM}};
  r_939_0 = _RAND_4438[0:0];
  _RAND_4439 = {1{`RANDOM}};
  r_939_1 = _RAND_4439[0:0];
  _RAND_4440 = {1{`RANDOM}};
  r_940_0 = _RAND_4440[0:0];
  _RAND_4441 = {1{`RANDOM}};
  r_940_1 = _RAND_4441[0:0];
  _RAND_4442 = {1{`RANDOM}};
  r_941_0 = _RAND_4442[0:0];
  _RAND_4443 = {1{`RANDOM}};
  r_941_1 = _RAND_4443[0:0];
  _RAND_4444 = {1{`RANDOM}};
  r_942_0 = _RAND_4444[0:0];
  _RAND_4445 = {1{`RANDOM}};
  r_942_1 = _RAND_4445[0:0];
  _RAND_4446 = {1{`RANDOM}};
  r_943_0 = _RAND_4446[0:0];
  _RAND_4447 = {1{`RANDOM}};
  r_943_1 = _RAND_4447[0:0];
  _RAND_4448 = {1{`RANDOM}};
  r_944_0 = _RAND_4448[0:0];
  _RAND_4449 = {1{`RANDOM}};
  r_944_1 = _RAND_4449[0:0];
  _RAND_4450 = {1{`RANDOM}};
  r_945_0 = _RAND_4450[0:0];
  _RAND_4451 = {1{`RANDOM}};
  r_945_1 = _RAND_4451[0:0];
  _RAND_4452 = {1{`RANDOM}};
  r_946_0 = _RAND_4452[0:0];
  _RAND_4453 = {1{`RANDOM}};
  r_946_1 = _RAND_4453[0:0];
  _RAND_4454 = {1{`RANDOM}};
  r_947_0 = _RAND_4454[0:0];
  _RAND_4455 = {1{`RANDOM}};
  r_947_1 = _RAND_4455[0:0];
  _RAND_4456 = {1{`RANDOM}};
  r_948_0 = _RAND_4456[0:0];
  _RAND_4457 = {1{`RANDOM}};
  r_948_1 = _RAND_4457[0:0];
  _RAND_4458 = {1{`RANDOM}};
  r_949_0 = _RAND_4458[0:0];
  _RAND_4459 = {1{`RANDOM}};
  r_949_1 = _RAND_4459[0:0];
  _RAND_4460 = {1{`RANDOM}};
  r_950_0 = _RAND_4460[0:0];
  _RAND_4461 = {1{`RANDOM}};
  r_950_1 = _RAND_4461[0:0];
  _RAND_4462 = {1{`RANDOM}};
  r_951_0 = _RAND_4462[0:0];
  _RAND_4463 = {1{`RANDOM}};
  r_951_1 = _RAND_4463[0:0];
  _RAND_4464 = {1{`RANDOM}};
  r_952_0 = _RAND_4464[0:0];
  _RAND_4465 = {1{`RANDOM}};
  r_952_1 = _RAND_4465[0:0];
  _RAND_4466 = {1{`RANDOM}};
  r_953_0 = _RAND_4466[0:0];
  _RAND_4467 = {1{`RANDOM}};
  r_953_1 = _RAND_4467[0:0];
  _RAND_4468 = {1{`RANDOM}};
  r_954_0 = _RAND_4468[0:0];
  _RAND_4469 = {1{`RANDOM}};
  r_954_1 = _RAND_4469[0:0];
  _RAND_4470 = {1{`RANDOM}};
  r_955_0 = _RAND_4470[0:0];
  _RAND_4471 = {1{`RANDOM}};
  r_955_1 = _RAND_4471[0:0];
  _RAND_4472 = {1{`RANDOM}};
  r_956_0 = _RAND_4472[0:0];
  _RAND_4473 = {1{`RANDOM}};
  r_956_1 = _RAND_4473[0:0];
  _RAND_4474 = {1{`RANDOM}};
  r_957_0 = _RAND_4474[0:0];
  _RAND_4475 = {1{`RANDOM}};
  r_957_1 = _RAND_4475[0:0];
  _RAND_4476 = {1{`RANDOM}};
  r_958_0 = _RAND_4476[0:0];
  _RAND_4477 = {1{`RANDOM}};
  r_958_1 = _RAND_4477[0:0];
  _RAND_4478 = {1{`RANDOM}};
  r_959_0 = _RAND_4478[0:0];
  _RAND_4479 = {1{`RANDOM}};
  r_959_1 = _RAND_4479[0:0];
  _RAND_4480 = {1{`RANDOM}};
  r_960_0 = _RAND_4480[0:0];
  _RAND_4481 = {1{`RANDOM}};
  r_960_1 = _RAND_4481[0:0];
  _RAND_4482 = {1{`RANDOM}};
  r_961_0 = _RAND_4482[0:0];
  _RAND_4483 = {1{`RANDOM}};
  r_961_1 = _RAND_4483[0:0];
  _RAND_4484 = {1{`RANDOM}};
  r_962_0 = _RAND_4484[0:0];
  _RAND_4485 = {1{`RANDOM}};
  r_962_1 = _RAND_4485[0:0];
  _RAND_4486 = {1{`RANDOM}};
  r_963_0 = _RAND_4486[0:0];
  _RAND_4487 = {1{`RANDOM}};
  r_963_1 = _RAND_4487[0:0];
  _RAND_4488 = {1{`RANDOM}};
  r_964_0 = _RAND_4488[0:0];
  _RAND_4489 = {1{`RANDOM}};
  r_964_1 = _RAND_4489[0:0];
  _RAND_4490 = {1{`RANDOM}};
  r_965_0 = _RAND_4490[0:0];
  _RAND_4491 = {1{`RANDOM}};
  r_965_1 = _RAND_4491[0:0];
  _RAND_4492 = {1{`RANDOM}};
  r_966_0 = _RAND_4492[0:0];
  _RAND_4493 = {1{`RANDOM}};
  r_966_1 = _RAND_4493[0:0];
  _RAND_4494 = {1{`RANDOM}};
  r_967_0 = _RAND_4494[0:0];
  _RAND_4495 = {1{`RANDOM}};
  r_967_1 = _RAND_4495[0:0];
  _RAND_4496 = {1{`RANDOM}};
  r_968_0 = _RAND_4496[0:0];
  _RAND_4497 = {1{`RANDOM}};
  r_968_1 = _RAND_4497[0:0];
  _RAND_4498 = {1{`RANDOM}};
  r_969_0 = _RAND_4498[0:0];
  _RAND_4499 = {1{`RANDOM}};
  r_969_1 = _RAND_4499[0:0];
  _RAND_4500 = {1{`RANDOM}};
  r_970_0 = _RAND_4500[0:0];
  _RAND_4501 = {1{`RANDOM}};
  r_970_1 = _RAND_4501[0:0];
  _RAND_4502 = {1{`RANDOM}};
  r_971_0 = _RAND_4502[0:0];
  _RAND_4503 = {1{`RANDOM}};
  r_971_1 = _RAND_4503[0:0];
  _RAND_4504 = {1{`RANDOM}};
  r_972_0 = _RAND_4504[0:0];
  _RAND_4505 = {1{`RANDOM}};
  r_972_1 = _RAND_4505[0:0];
  _RAND_4506 = {1{`RANDOM}};
  r_973_0 = _RAND_4506[0:0];
  _RAND_4507 = {1{`RANDOM}};
  r_973_1 = _RAND_4507[0:0];
  _RAND_4508 = {1{`RANDOM}};
  r_974_0 = _RAND_4508[0:0];
  _RAND_4509 = {1{`RANDOM}};
  r_974_1 = _RAND_4509[0:0];
  _RAND_4510 = {1{`RANDOM}};
  r_975_0 = _RAND_4510[0:0];
  _RAND_4511 = {1{`RANDOM}};
  r_975_1 = _RAND_4511[0:0];
  _RAND_4512 = {1{`RANDOM}};
  r_976_0 = _RAND_4512[0:0];
  _RAND_4513 = {1{`RANDOM}};
  r_976_1 = _RAND_4513[0:0];
  _RAND_4514 = {1{`RANDOM}};
  r_977_0 = _RAND_4514[0:0];
  _RAND_4515 = {1{`RANDOM}};
  r_977_1 = _RAND_4515[0:0];
  _RAND_4516 = {1{`RANDOM}};
  r_978_0 = _RAND_4516[0:0];
  _RAND_4517 = {1{`RANDOM}};
  r_978_1 = _RAND_4517[0:0];
  _RAND_4518 = {1{`RANDOM}};
  r_979_0 = _RAND_4518[0:0];
  _RAND_4519 = {1{`RANDOM}};
  r_979_1 = _RAND_4519[0:0];
  _RAND_4520 = {1{`RANDOM}};
  r_980_0 = _RAND_4520[0:0];
  _RAND_4521 = {1{`RANDOM}};
  r_980_1 = _RAND_4521[0:0];
  _RAND_4522 = {1{`RANDOM}};
  r_981_0 = _RAND_4522[0:0];
  _RAND_4523 = {1{`RANDOM}};
  r_981_1 = _RAND_4523[0:0];
  _RAND_4524 = {1{`RANDOM}};
  r_982_0 = _RAND_4524[0:0];
  _RAND_4525 = {1{`RANDOM}};
  r_982_1 = _RAND_4525[0:0];
  _RAND_4526 = {1{`RANDOM}};
  r_983_0 = _RAND_4526[0:0];
  _RAND_4527 = {1{`RANDOM}};
  r_983_1 = _RAND_4527[0:0];
  _RAND_4528 = {1{`RANDOM}};
  r_984_0 = _RAND_4528[0:0];
  _RAND_4529 = {1{`RANDOM}};
  r_984_1 = _RAND_4529[0:0];
  _RAND_4530 = {1{`RANDOM}};
  r_985_0 = _RAND_4530[0:0];
  _RAND_4531 = {1{`RANDOM}};
  r_985_1 = _RAND_4531[0:0];
  _RAND_4532 = {1{`RANDOM}};
  r_986_0 = _RAND_4532[0:0];
  _RAND_4533 = {1{`RANDOM}};
  r_986_1 = _RAND_4533[0:0];
  _RAND_4534 = {1{`RANDOM}};
  r_987_0 = _RAND_4534[0:0];
  _RAND_4535 = {1{`RANDOM}};
  r_987_1 = _RAND_4535[0:0];
  _RAND_4536 = {1{`RANDOM}};
  r_988_0 = _RAND_4536[0:0];
  _RAND_4537 = {1{`RANDOM}};
  r_988_1 = _RAND_4537[0:0];
  _RAND_4538 = {1{`RANDOM}};
  r_989_0 = _RAND_4538[0:0];
  _RAND_4539 = {1{`RANDOM}};
  r_989_1 = _RAND_4539[0:0];
  _RAND_4540 = {1{`RANDOM}};
  r_990_0 = _RAND_4540[0:0];
  _RAND_4541 = {1{`RANDOM}};
  r_990_1 = _RAND_4541[0:0];
  _RAND_4542 = {1{`RANDOM}};
  r_991_0 = _RAND_4542[0:0];
  _RAND_4543 = {1{`RANDOM}};
  r_991_1 = _RAND_4543[0:0];
  _RAND_4544 = {1{`RANDOM}};
  r_992_0 = _RAND_4544[0:0];
  _RAND_4545 = {1{`RANDOM}};
  r_992_1 = _RAND_4545[0:0];
  _RAND_4546 = {1{`RANDOM}};
  r_993_0 = _RAND_4546[0:0];
  _RAND_4547 = {1{`RANDOM}};
  r_993_1 = _RAND_4547[0:0];
  _RAND_4548 = {1{`RANDOM}};
  r_994_0 = _RAND_4548[0:0];
  _RAND_4549 = {1{`RANDOM}};
  r_994_1 = _RAND_4549[0:0];
  _RAND_4550 = {1{`RANDOM}};
  r_995_0 = _RAND_4550[0:0];
  _RAND_4551 = {1{`RANDOM}};
  r_995_1 = _RAND_4551[0:0];
  _RAND_4552 = {1{`RANDOM}};
  r_996_0 = _RAND_4552[0:0];
  _RAND_4553 = {1{`RANDOM}};
  r_996_1 = _RAND_4553[0:0];
  _RAND_4554 = {1{`RANDOM}};
  r_997_0 = _RAND_4554[0:0];
  _RAND_4555 = {1{`RANDOM}};
  r_997_1 = _RAND_4555[0:0];
  _RAND_4556 = {1{`RANDOM}};
  r_998_0 = _RAND_4556[0:0];
  _RAND_4557 = {1{`RANDOM}};
  r_998_1 = _RAND_4557[0:0];
  _RAND_4558 = {1{`RANDOM}};
  r_999_0 = _RAND_4558[0:0];
  _RAND_4559 = {1{`RANDOM}};
  r_999_1 = _RAND_4559[0:0];
  _RAND_4560 = {1{`RANDOM}};
  r_1000_0 = _RAND_4560[0:0];
  _RAND_4561 = {1{`RANDOM}};
  r_1000_1 = _RAND_4561[0:0];
  _RAND_4562 = {1{`RANDOM}};
  r_1001_0 = _RAND_4562[0:0];
  _RAND_4563 = {1{`RANDOM}};
  r_1001_1 = _RAND_4563[0:0];
  _RAND_4564 = {1{`RANDOM}};
  r_1002_0 = _RAND_4564[0:0];
  _RAND_4565 = {1{`RANDOM}};
  r_1002_1 = _RAND_4565[0:0];
  _RAND_4566 = {1{`RANDOM}};
  r_1003_0 = _RAND_4566[0:0];
  _RAND_4567 = {1{`RANDOM}};
  r_1003_1 = _RAND_4567[0:0];
  _RAND_4568 = {1{`RANDOM}};
  r_1004_0 = _RAND_4568[0:0];
  _RAND_4569 = {1{`RANDOM}};
  r_1004_1 = _RAND_4569[0:0];
  _RAND_4570 = {1{`RANDOM}};
  r_1005_0 = _RAND_4570[0:0];
  _RAND_4571 = {1{`RANDOM}};
  r_1005_1 = _RAND_4571[0:0];
  _RAND_4572 = {1{`RANDOM}};
  r_1006_0 = _RAND_4572[0:0];
  _RAND_4573 = {1{`RANDOM}};
  r_1006_1 = _RAND_4573[0:0];
  _RAND_4574 = {1{`RANDOM}};
  r_1007_0 = _RAND_4574[0:0];
  _RAND_4575 = {1{`RANDOM}};
  r_1007_1 = _RAND_4575[0:0];
  _RAND_4576 = {1{`RANDOM}};
  r_1008_0 = _RAND_4576[0:0];
  _RAND_4577 = {1{`RANDOM}};
  r_1008_1 = _RAND_4577[0:0];
  _RAND_4578 = {1{`RANDOM}};
  r_1009_0 = _RAND_4578[0:0];
  _RAND_4579 = {1{`RANDOM}};
  r_1009_1 = _RAND_4579[0:0];
  _RAND_4580 = {1{`RANDOM}};
  r_1010_0 = _RAND_4580[0:0];
  _RAND_4581 = {1{`RANDOM}};
  r_1010_1 = _RAND_4581[0:0];
  _RAND_4582 = {1{`RANDOM}};
  r_1011_0 = _RAND_4582[0:0];
  _RAND_4583 = {1{`RANDOM}};
  r_1011_1 = _RAND_4583[0:0];
  _RAND_4584 = {1{`RANDOM}};
  r_1012_0 = _RAND_4584[0:0];
  _RAND_4585 = {1{`RANDOM}};
  r_1012_1 = _RAND_4585[0:0];
  _RAND_4586 = {1{`RANDOM}};
  r_1013_0 = _RAND_4586[0:0];
  _RAND_4587 = {1{`RANDOM}};
  r_1013_1 = _RAND_4587[0:0];
  _RAND_4588 = {1{`RANDOM}};
  r_1014_0 = _RAND_4588[0:0];
  _RAND_4589 = {1{`RANDOM}};
  r_1014_1 = _RAND_4589[0:0];
  _RAND_4590 = {1{`RANDOM}};
  r_1015_0 = _RAND_4590[0:0];
  _RAND_4591 = {1{`RANDOM}};
  r_1015_1 = _RAND_4591[0:0];
  _RAND_4592 = {1{`RANDOM}};
  r_1016_0 = _RAND_4592[0:0];
  _RAND_4593 = {1{`RANDOM}};
  r_1016_1 = _RAND_4593[0:0];
  _RAND_4594 = {1{`RANDOM}};
  r_1017_0 = _RAND_4594[0:0];
  _RAND_4595 = {1{`RANDOM}};
  r_1017_1 = _RAND_4595[0:0];
  _RAND_4596 = {1{`RANDOM}};
  r_1018_0 = _RAND_4596[0:0];
  _RAND_4597 = {1{`RANDOM}};
  r_1018_1 = _RAND_4597[0:0];
  _RAND_4598 = {1{`RANDOM}};
  r_1019_0 = _RAND_4598[0:0];
  _RAND_4599 = {1{`RANDOM}};
  r_1019_1 = _RAND_4599[0:0];
  _RAND_4600 = {1{`RANDOM}};
  r_1020_0 = _RAND_4600[0:0];
  _RAND_4601 = {1{`RANDOM}};
  r_1020_1 = _RAND_4601[0:0];
  _RAND_4602 = {1{`RANDOM}};
  r_1021_0 = _RAND_4602[0:0];
  _RAND_4603 = {1{`RANDOM}};
  r_1021_1 = _RAND_4603[0:0];
  _RAND_4604 = {1{`RANDOM}};
  r_1022_0 = _RAND_4604[0:0];
  _RAND_4605 = {1{`RANDOM}};
  r_1022_1 = _RAND_4605[0:0];
  _RAND_4606 = {1{`RANDOM}};
  r_1023_0 = _RAND_4606[0:0];
  _RAND_4607 = {1{`RANDOM}};
  r_1023_1 = _RAND_4607[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module gemmini(
  input         clock,
  input         reset,
  input  [7:0]  io_in_a_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_a_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_b_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [7:0]  io_in_d_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_0_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_0_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_0_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_0_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_0_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_0_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_1_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_1_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_1_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_1_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_1_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_1_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_2_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_2_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_2_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_2_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_2_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_2_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_3_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_3_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_3_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_3_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_3_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_3_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_4_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_4_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_4_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_4_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_4_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_4_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_5_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_5_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_5_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_5_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_5_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_5_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_6_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_6_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_6_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_6_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_6_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_6_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_7_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_7_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_7_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_7_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_7_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_7_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_8_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_8_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_8_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_8_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_8_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_8_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_9_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_9_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_9_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_9_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_9_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_9_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_10_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_10_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_10_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_10_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_10_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_10_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_11_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_11_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_11_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_11_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_11_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_11_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_12_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_12_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_12_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_12_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_12_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_12_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_13_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_13_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_13_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_13_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_13_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_13_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_14_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_14_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_14_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_14_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_14_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_14_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_15_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_15_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_15_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_15_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_control_15_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [4:0]  io_in_control_15_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input  [1:0]  io_in_id_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_last_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  input         io_in_valid_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_b_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [19:0] io_out_c_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_valid_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_0_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_0_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_0_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_0_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_0_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_0_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_1_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_1_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_1_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_1_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_1_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_1_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_2_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_2_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_2_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_2_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_2_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_2_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_3_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_3_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_3_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_3_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_3_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_3_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_4_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_4_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_4_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_4_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_4_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_4_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_5_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_5_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_5_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_5_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_5_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_5_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_6_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_6_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_6_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_6_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_6_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_6_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_7_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_7_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_7_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_7_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_7_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_7_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_8_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_8_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_8_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_8_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_8_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_8_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_9_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_9_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_9_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_9_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_9_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_9_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_10_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_10_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_10_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_10_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_10_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_10_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_11_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_11_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_11_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_11_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_11_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_11_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_12_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_12_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_12_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_12_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_12_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_12_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_13_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_13_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_13_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_13_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_13_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_13_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_14_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_14_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_14_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_14_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_14_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_14_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_15_0_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_15_0_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_15_0_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_15_1_dataflow, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_control_15_1_propagate, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [4:0]  io_out_control_15_1_shift, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output [1:0]  io_out_id_15_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_0_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_0_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_1_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_1_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_2_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_2_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_3_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_3_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_4_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_4_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_5_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_5_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_6_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_6_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_7_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_7_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_8_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_8_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_9_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_9_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_10_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_10_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_11_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_11_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_12_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_12_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_13_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_13_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_14_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_14_1, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_15_0, // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
  output        io_out_last_15_1 // @[src/main/scala/gemmini/GemminiMeshTop.scala 42:14]
);
  wire  mesh_clock; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_a_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_b_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [7:0] mesh_io_in_d_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_0_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_0_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_0_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_0_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_0_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_0_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_1_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_1_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_1_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_1_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_1_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_1_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_2_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_2_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_2_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_2_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_2_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_2_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_3_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_3_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_3_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_3_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_3_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_3_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_4_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_4_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_4_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_4_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_4_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_4_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_5_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_5_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_5_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_5_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_5_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_5_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_6_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_6_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_6_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_6_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_6_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_6_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_7_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_7_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_7_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_7_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_7_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_7_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_8_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_8_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_8_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_8_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_8_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_8_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_9_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_9_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_9_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_9_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_9_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_9_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_10_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_10_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_10_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_10_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_10_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_10_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_11_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_11_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_11_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_11_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_11_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_11_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_12_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_12_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_12_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_12_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_12_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_12_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_13_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_13_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_13_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_13_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_13_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_13_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_14_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_14_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_14_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_14_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_14_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_14_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_15_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_15_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_15_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_15_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_control_15_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_in_control_15_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_in_id_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_last_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_b_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [19:0] mesh_io_out_c_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_in_valid_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_valid_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_0_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_0_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_0_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_0_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_0_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_0_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_1_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_1_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_1_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_1_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_1_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_1_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_2_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_2_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_2_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_2_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_2_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_2_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_3_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_3_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_3_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_3_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_3_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_3_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_4_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_4_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_4_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_4_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_4_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_4_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_5_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_5_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_5_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_5_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_5_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_5_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_6_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_6_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_6_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_6_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_6_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_6_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_7_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_7_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_7_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_7_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_7_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_7_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_8_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_8_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_8_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_8_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_8_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_8_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_9_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_9_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_9_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_9_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_9_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_9_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_10_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_10_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_10_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_10_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_10_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_10_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_11_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_11_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_11_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_11_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_11_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_11_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_12_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_12_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_12_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_12_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_12_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_12_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_13_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_13_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_13_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_13_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_13_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_13_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_14_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_14_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_14_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_14_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_14_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_14_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_15_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_15_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_15_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_15_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_control_15_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [4:0] mesh_io_out_control_15_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire [1:0] mesh_io_out_id_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  wire  mesh_io_out_last_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
  Mesh mesh ( // @[src/main/scala/gemmini/GemminiMeshTop.scala 26:20]
    .clock(mesh_clock),
    .io_in_a_0_0(mesh_io_in_a_0_0),
    .io_in_a_0_1(mesh_io_in_a_0_1),
    .io_in_a_1_0(mesh_io_in_a_1_0),
    .io_in_a_1_1(mesh_io_in_a_1_1),
    .io_in_a_2_0(mesh_io_in_a_2_0),
    .io_in_a_2_1(mesh_io_in_a_2_1),
    .io_in_a_3_0(mesh_io_in_a_3_0),
    .io_in_a_3_1(mesh_io_in_a_3_1),
    .io_in_a_4_0(mesh_io_in_a_4_0),
    .io_in_a_4_1(mesh_io_in_a_4_1),
    .io_in_a_5_0(mesh_io_in_a_5_0),
    .io_in_a_5_1(mesh_io_in_a_5_1),
    .io_in_a_6_0(mesh_io_in_a_6_0),
    .io_in_a_6_1(mesh_io_in_a_6_1),
    .io_in_a_7_0(mesh_io_in_a_7_0),
    .io_in_a_7_1(mesh_io_in_a_7_1),
    .io_in_a_8_0(mesh_io_in_a_8_0),
    .io_in_a_8_1(mesh_io_in_a_8_1),
    .io_in_a_9_0(mesh_io_in_a_9_0),
    .io_in_a_9_1(mesh_io_in_a_9_1),
    .io_in_a_10_0(mesh_io_in_a_10_0),
    .io_in_a_10_1(mesh_io_in_a_10_1),
    .io_in_a_11_0(mesh_io_in_a_11_0),
    .io_in_a_11_1(mesh_io_in_a_11_1),
    .io_in_a_12_0(mesh_io_in_a_12_0),
    .io_in_a_12_1(mesh_io_in_a_12_1),
    .io_in_a_13_0(mesh_io_in_a_13_0),
    .io_in_a_13_1(mesh_io_in_a_13_1),
    .io_in_a_14_0(mesh_io_in_a_14_0),
    .io_in_a_14_1(mesh_io_in_a_14_1),
    .io_in_a_15_0(mesh_io_in_a_15_0),
    .io_in_a_15_1(mesh_io_in_a_15_1),
    .io_in_b_0_0(mesh_io_in_b_0_0),
    .io_in_b_0_1(mesh_io_in_b_0_1),
    .io_in_b_1_0(mesh_io_in_b_1_0),
    .io_in_b_1_1(mesh_io_in_b_1_1),
    .io_in_b_2_0(mesh_io_in_b_2_0),
    .io_in_b_2_1(mesh_io_in_b_2_1),
    .io_in_b_3_0(mesh_io_in_b_3_0),
    .io_in_b_3_1(mesh_io_in_b_3_1),
    .io_in_b_4_0(mesh_io_in_b_4_0),
    .io_in_b_4_1(mesh_io_in_b_4_1),
    .io_in_b_5_0(mesh_io_in_b_5_0),
    .io_in_b_5_1(mesh_io_in_b_5_1),
    .io_in_b_6_0(mesh_io_in_b_6_0),
    .io_in_b_6_1(mesh_io_in_b_6_1),
    .io_in_b_7_0(mesh_io_in_b_7_0),
    .io_in_b_7_1(mesh_io_in_b_7_1),
    .io_in_b_8_0(mesh_io_in_b_8_0),
    .io_in_b_8_1(mesh_io_in_b_8_1),
    .io_in_b_9_0(mesh_io_in_b_9_0),
    .io_in_b_9_1(mesh_io_in_b_9_1),
    .io_in_b_10_0(mesh_io_in_b_10_0),
    .io_in_b_10_1(mesh_io_in_b_10_1),
    .io_in_b_11_0(mesh_io_in_b_11_0),
    .io_in_b_11_1(mesh_io_in_b_11_1),
    .io_in_b_12_0(mesh_io_in_b_12_0),
    .io_in_b_12_1(mesh_io_in_b_12_1),
    .io_in_b_13_0(mesh_io_in_b_13_0),
    .io_in_b_13_1(mesh_io_in_b_13_1),
    .io_in_b_14_0(mesh_io_in_b_14_0),
    .io_in_b_14_1(mesh_io_in_b_14_1),
    .io_in_b_15_0(mesh_io_in_b_15_0),
    .io_in_b_15_1(mesh_io_in_b_15_1),
    .io_in_d_0_0(mesh_io_in_d_0_0),
    .io_in_d_0_1(mesh_io_in_d_0_1),
    .io_in_d_1_0(mesh_io_in_d_1_0),
    .io_in_d_1_1(mesh_io_in_d_1_1),
    .io_in_d_2_0(mesh_io_in_d_2_0),
    .io_in_d_2_1(mesh_io_in_d_2_1),
    .io_in_d_3_0(mesh_io_in_d_3_0),
    .io_in_d_3_1(mesh_io_in_d_3_1),
    .io_in_d_4_0(mesh_io_in_d_4_0),
    .io_in_d_4_1(mesh_io_in_d_4_1),
    .io_in_d_5_0(mesh_io_in_d_5_0),
    .io_in_d_5_1(mesh_io_in_d_5_1),
    .io_in_d_6_0(mesh_io_in_d_6_0),
    .io_in_d_6_1(mesh_io_in_d_6_1),
    .io_in_d_7_0(mesh_io_in_d_7_0),
    .io_in_d_7_1(mesh_io_in_d_7_1),
    .io_in_d_8_0(mesh_io_in_d_8_0),
    .io_in_d_8_1(mesh_io_in_d_8_1),
    .io_in_d_9_0(mesh_io_in_d_9_0),
    .io_in_d_9_1(mesh_io_in_d_9_1),
    .io_in_d_10_0(mesh_io_in_d_10_0),
    .io_in_d_10_1(mesh_io_in_d_10_1),
    .io_in_d_11_0(mesh_io_in_d_11_0),
    .io_in_d_11_1(mesh_io_in_d_11_1),
    .io_in_d_12_0(mesh_io_in_d_12_0),
    .io_in_d_12_1(mesh_io_in_d_12_1),
    .io_in_d_13_0(mesh_io_in_d_13_0),
    .io_in_d_13_1(mesh_io_in_d_13_1),
    .io_in_d_14_0(mesh_io_in_d_14_0),
    .io_in_d_14_1(mesh_io_in_d_14_1),
    .io_in_d_15_0(mesh_io_in_d_15_0),
    .io_in_d_15_1(mesh_io_in_d_15_1),
    .io_in_control_0_0_dataflow(mesh_io_in_control_0_0_dataflow),
    .io_in_control_0_0_propagate(mesh_io_in_control_0_0_propagate),
    .io_in_control_0_0_shift(mesh_io_in_control_0_0_shift),
    .io_in_control_0_1_dataflow(mesh_io_in_control_0_1_dataflow),
    .io_in_control_0_1_propagate(mesh_io_in_control_0_1_propagate),
    .io_in_control_0_1_shift(mesh_io_in_control_0_1_shift),
    .io_in_control_1_0_dataflow(mesh_io_in_control_1_0_dataflow),
    .io_in_control_1_0_propagate(mesh_io_in_control_1_0_propagate),
    .io_in_control_1_0_shift(mesh_io_in_control_1_0_shift),
    .io_in_control_1_1_dataflow(mesh_io_in_control_1_1_dataflow),
    .io_in_control_1_1_propagate(mesh_io_in_control_1_1_propagate),
    .io_in_control_1_1_shift(mesh_io_in_control_1_1_shift),
    .io_in_control_2_0_dataflow(mesh_io_in_control_2_0_dataflow),
    .io_in_control_2_0_propagate(mesh_io_in_control_2_0_propagate),
    .io_in_control_2_0_shift(mesh_io_in_control_2_0_shift),
    .io_in_control_2_1_dataflow(mesh_io_in_control_2_1_dataflow),
    .io_in_control_2_1_propagate(mesh_io_in_control_2_1_propagate),
    .io_in_control_2_1_shift(mesh_io_in_control_2_1_shift),
    .io_in_control_3_0_dataflow(mesh_io_in_control_3_0_dataflow),
    .io_in_control_3_0_propagate(mesh_io_in_control_3_0_propagate),
    .io_in_control_3_0_shift(mesh_io_in_control_3_0_shift),
    .io_in_control_3_1_dataflow(mesh_io_in_control_3_1_dataflow),
    .io_in_control_3_1_propagate(mesh_io_in_control_3_1_propagate),
    .io_in_control_3_1_shift(mesh_io_in_control_3_1_shift),
    .io_in_control_4_0_dataflow(mesh_io_in_control_4_0_dataflow),
    .io_in_control_4_0_propagate(mesh_io_in_control_4_0_propagate),
    .io_in_control_4_0_shift(mesh_io_in_control_4_0_shift),
    .io_in_control_4_1_dataflow(mesh_io_in_control_4_1_dataflow),
    .io_in_control_4_1_propagate(mesh_io_in_control_4_1_propagate),
    .io_in_control_4_1_shift(mesh_io_in_control_4_1_shift),
    .io_in_control_5_0_dataflow(mesh_io_in_control_5_0_dataflow),
    .io_in_control_5_0_propagate(mesh_io_in_control_5_0_propagate),
    .io_in_control_5_0_shift(mesh_io_in_control_5_0_shift),
    .io_in_control_5_1_dataflow(mesh_io_in_control_5_1_dataflow),
    .io_in_control_5_1_propagate(mesh_io_in_control_5_1_propagate),
    .io_in_control_5_1_shift(mesh_io_in_control_5_1_shift),
    .io_in_control_6_0_dataflow(mesh_io_in_control_6_0_dataflow),
    .io_in_control_6_0_propagate(mesh_io_in_control_6_0_propagate),
    .io_in_control_6_0_shift(mesh_io_in_control_6_0_shift),
    .io_in_control_6_1_dataflow(mesh_io_in_control_6_1_dataflow),
    .io_in_control_6_1_propagate(mesh_io_in_control_6_1_propagate),
    .io_in_control_6_1_shift(mesh_io_in_control_6_1_shift),
    .io_in_control_7_0_dataflow(mesh_io_in_control_7_0_dataflow),
    .io_in_control_7_0_propagate(mesh_io_in_control_7_0_propagate),
    .io_in_control_7_0_shift(mesh_io_in_control_7_0_shift),
    .io_in_control_7_1_dataflow(mesh_io_in_control_7_1_dataflow),
    .io_in_control_7_1_propagate(mesh_io_in_control_7_1_propagate),
    .io_in_control_7_1_shift(mesh_io_in_control_7_1_shift),
    .io_in_control_8_0_dataflow(mesh_io_in_control_8_0_dataflow),
    .io_in_control_8_0_propagate(mesh_io_in_control_8_0_propagate),
    .io_in_control_8_0_shift(mesh_io_in_control_8_0_shift),
    .io_in_control_8_1_dataflow(mesh_io_in_control_8_1_dataflow),
    .io_in_control_8_1_propagate(mesh_io_in_control_8_1_propagate),
    .io_in_control_8_1_shift(mesh_io_in_control_8_1_shift),
    .io_in_control_9_0_dataflow(mesh_io_in_control_9_0_dataflow),
    .io_in_control_9_0_propagate(mesh_io_in_control_9_0_propagate),
    .io_in_control_9_0_shift(mesh_io_in_control_9_0_shift),
    .io_in_control_9_1_dataflow(mesh_io_in_control_9_1_dataflow),
    .io_in_control_9_1_propagate(mesh_io_in_control_9_1_propagate),
    .io_in_control_9_1_shift(mesh_io_in_control_9_1_shift),
    .io_in_control_10_0_dataflow(mesh_io_in_control_10_0_dataflow),
    .io_in_control_10_0_propagate(mesh_io_in_control_10_0_propagate),
    .io_in_control_10_0_shift(mesh_io_in_control_10_0_shift),
    .io_in_control_10_1_dataflow(mesh_io_in_control_10_1_dataflow),
    .io_in_control_10_1_propagate(mesh_io_in_control_10_1_propagate),
    .io_in_control_10_1_shift(mesh_io_in_control_10_1_shift),
    .io_in_control_11_0_dataflow(mesh_io_in_control_11_0_dataflow),
    .io_in_control_11_0_propagate(mesh_io_in_control_11_0_propagate),
    .io_in_control_11_0_shift(mesh_io_in_control_11_0_shift),
    .io_in_control_11_1_dataflow(mesh_io_in_control_11_1_dataflow),
    .io_in_control_11_1_propagate(mesh_io_in_control_11_1_propagate),
    .io_in_control_11_1_shift(mesh_io_in_control_11_1_shift),
    .io_in_control_12_0_dataflow(mesh_io_in_control_12_0_dataflow),
    .io_in_control_12_0_propagate(mesh_io_in_control_12_0_propagate),
    .io_in_control_12_0_shift(mesh_io_in_control_12_0_shift),
    .io_in_control_12_1_dataflow(mesh_io_in_control_12_1_dataflow),
    .io_in_control_12_1_propagate(mesh_io_in_control_12_1_propagate),
    .io_in_control_12_1_shift(mesh_io_in_control_12_1_shift),
    .io_in_control_13_0_dataflow(mesh_io_in_control_13_0_dataflow),
    .io_in_control_13_0_propagate(mesh_io_in_control_13_0_propagate),
    .io_in_control_13_0_shift(mesh_io_in_control_13_0_shift),
    .io_in_control_13_1_dataflow(mesh_io_in_control_13_1_dataflow),
    .io_in_control_13_1_propagate(mesh_io_in_control_13_1_propagate),
    .io_in_control_13_1_shift(mesh_io_in_control_13_1_shift),
    .io_in_control_14_0_dataflow(mesh_io_in_control_14_0_dataflow),
    .io_in_control_14_0_propagate(mesh_io_in_control_14_0_propagate),
    .io_in_control_14_0_shift(mesh_io_in_control_14_0_shift),
    .io_in_control_14_1_dataflow(mesh_io_in_control_14_1_dataflow),
    .io_in_control_14_1_propagate(mesh_io_in_control_14_1_propagate),
    .io_in_control_14_1_shift(mesh_io_in_control_14_1_shift),
    .io_in_control_15_0_dataflow(mesh_io_in_control_15_0_dataflow),
    .io_in_control_15_0_propagate(mesh_io_in_control_15_0_propagate),
    .io_in_control_15_0_shift(mesh_io_in_control_15_0_shift),
    .io_in_control_15_1_dataflow(mesh_io_in_control_15_1_dataflow),
    .io_in_control_15_1_propagate(mesh_io_in_control_15_1_propagate),
    .io_in_control_15_1_shift(mesh_io_in_control_15_1_shift),
    .io_in_id_0_0(mesh_io_in_id_0_0),
    .io_in_id_0_1(mesh_io_in_id_0_1),
    .io_in_id_1_0(mesh_io_in_id_1_0),
    .io_in_id_1_1(mesh_io_in_id_1_1),
    .io_in_id_2_0(mesh_io_in_id_2_0),
    .io_in_id_2_1(mesh_io_in_id_2_1),
    .io_in_id_3_0(mesh_io_in_id_3_0),
    .io_in_id_3_1(mesh_io_in_id_3_1),
    .io_in_id_4_0(mesh_io_in_id_4_0),
    .io_in_id_4_1(mesh_io_in_id_4_1),
    .io_in_id_5_0(mesh_io_in_id_5_0),
    .io_in_id_5_1(mesh_io_in_id_5_1),
    .io_in_id_6_0(mesh_io_in_id_6_0),
    .io_in_id_6_1(mesh_io_in_id_6_1),
    .io_in_id_7_0(mesh_io_in_id_7_0),
    .io_in_id_7_1(mesh_io_in_id_7_1),
    .io_in_id_8_0(mesh_io_in_id_8_0),
    .io_in_id_8_1(mesh_io_in_id_8_1),
    .io_in_id_9_0(mesh_io_in_id_9_0),
    .io_in_id_9_1(mesh_io_in_id_9_1),
    .io_in_id_10_0(mesh_io_in_id_10_0),
    .io_in_id_10_1(mesh_io_in_id_10_1),
    .io_in_id_11_0(mesh_io_in_id_11_0),
    .io_in_id_11_1(mesh_io_in_id_11_1),
    .io_in_id_12_0(mesh_io_in_id_12_0),
    .io_in_id_12_1(mesh_io_in_id_12_1),
    .io_in_id_13_0(mesh_io_in_id_13_0),
    .io_in_id_13_1(mesh_io_in_id_13_1),
    .io_in_id_14_0(mesh_io_in_id_14_0),
    .io_in_id_14_1(mesh_io_in_id_14_1),
    .io_in_id_15_0(mesh_io_in_id_15_0),
    .io_in_id_15_1(mesh_io_in_id_15_1),
    .io_in_last_0_0(mesh_io_in_last_0_0),
    .io_in_last_0_1(mesh_io_in_last_0_1),
    .io_in_last_1_0(mesh_io_in_last_1_0),
    .io_in_last_1_1(mesh_io_in_last_1_1),
    .io_in_last_2_0(mesh_io_in_last_2_0),
    .io_in_last_2_1(mesh_io_in_last_2_1),
    .io_in_last_3_0(mesh_io_in_last_3_0),
    .io_in_last_3_1(mesh_io_in_last_3_1),
    .io_in_last_4_0(mesh_io_in_last_4_0),
    .io_in_last_4_1(mesh_io_in_last_4_1),
    .io_in_last_5_0(mesh_io_in_last_5_0),
    .io_in_last_5_1(mesh_io_in_last_5_1),
    .io_in_last_6_0(mesh_io_in_last_6_0),
    .io_in_last_6_1(mesh_io_in_last_6_1),
    .io_in_last_7_0(mesh_io_in_last_7_0),
    .io_in_last_7_1(mesh_io_in_last_7_1),
    .io_in_last_8_0(mesh_io_in_last_8_0),
    .io_in_last_8_1(mesh_io_in_last_8_1),
    .io_in_last_9_0(mesh_io_in_last_9_0),
    .io_in_last_9_1(mesh_io_in_last_9_1),
    .io_in_last_10_0(mesh_io_in_last_10_0),
    .io_in_last_10_1(mesh_io_in_last_10_1),
    .io_in_last_11_0(mesh_io_in_last_11_0),
    .io_in_last_11_1(mesh_io_in_last_11_1),
    .io_in_last_12_0(mesh_io_in_last_12_0),
    .io_in_last_12_1(mesh_io_in_last_12_1),
    .io_in_last_13_0(mesh_io_in_last_13_0),
    .io_in_last_13_1(mesh_io_in_last_13_1),
    .io_in_last_14_0(mesh_io_in_last_14_0),
    .io_in_last_14_1(mesh_io_in_last_14_1),
    .io_in_last_15_0(mesh_io_in_last_15_0),
    .io_in_last_15_1(mesh_io_in_last_15_1),
    .io_out_b_0_0(mesh_io_out_b_0_0),
    .io_out_b_0_1(mesh_io_out_b_0_1),
    .io_out_b_1_0(mesh_io_out_b_1_0),
    .io_out_b_1_1(mesh_io_out_b_1_1),
    .io_out_b_2_0(mesh_io_out_b_2_0),
    .io_out_b_2_1(mesh_io_out_b_2_1),
    .io_out_b_3_0(mesh_io_out_b_3_0),
    .io_out_b_3_1(mesh_io_out_b_3_1),
    .io_out_b_4_0(mesh_io_out_b_4_0),
    .io_out_b_4_1(mesh_io_out_b_4_1),
    .io_out_b_5_0(mesh_io_out_b_5_0),
    .io_out_b_5_1(mesh_io_out_b_5_1),
    .io_out_b_6_0(mesh_io_out_b_6_0),
    .io_out_b_6_1(mesh_io_out_b_6_1),
    .io_out_b_7_0(mesh_io_out_b_7_0),
    .io_out_b_7_1(mesh_io_out_b_7_1),
    .io_out_b_8_0(mesh_io_out_b_8_0),
    .io_out_b_8_1(mesh_io_out_b_8_1),
    .io_out_b_9_0(mesh_io_out_b_9_0),
    .io_out_b_9_1(mesh_io_out_b_9_1),
    .io_out_b_10_0(mesh_io_out_b_10_0),
    .io_out_b_10_1(mesh_io_out_b_10_1),
    .io_out_b_11_0(mesh_io_out_b_11_0),
    .io_out_b_11_1(mesh_io_out_b_11_1),
    .io_out_b_12_0(mesh_io_out_b_12_0),
    .io_out_b_12_1(mesh_io_out_b_12_1),
    .io_out_b_13_0(mesh_io_out_b_13_0),
    .io_out_b_13_1(mesh_io_out_b_13_1),
    .io_out_b_14_0(mesh_io_out_b_14_0),
    .io_out_b_14_1(mesh_io_out_b_14_1),
    .io_out_b_15_0(mesh_io_out_b_15_0),
    .io_out_b_15_1(mesh_io_out_b_15_1),
    .io_out_c_0_0(mesh_io_out_c_0_0),
    .io_out_c_0_1(mesh_io_out_c_0_1),
    .io_out_c_1_0(mesh_io_out_c_1_0),
    .io_out_c_1_1(mesh_io_out_c_1_1),
    .io_out_c_2_0(mesh_io_out_c_2_0),
    .io_out_c_2_1(mesh_io_out_c_2_1),
    .io_out_c_3_0(mesh_io_out_c_3_0),
    .io_out_c_3_1(mesh_io_out_c_3_1),
    .io_out_c_4_0(mesh_io_out_c_4_0),
    .io_out_c_4_1(mesh_io_out_c_4_1),
    .io_out_c_5_0(mesh_io_out_c_5_0),
    .io_out_c_5_1(mesh_io_out_c_5_1),
    .io_out_c_6_0(mesh_io_out_c_6_0),
    .io_out_c_6_1(mesh_io_out_c_6_1),
    .io_out_c_7_0(mesh_io_out_c_7_0),
    .io_out_c_7_1(mesh_io_out_c_7_1),
    .io_out_c_8_0(mesh_io_out_c_8_0),
    .io_out_c_8_1(mesh_io_out_c_8_1),
    .io_out_c_9_0(mesh_io_out_c_9_0),
    .io_out_c_9_1(mesh_io_out_c_9_1),
    .io_out_c_10_0(mesh_io_out_c_10_0),
    .io_out_c_10_1(mesh_io_out_c_10_1),
    .io_out_c_11_0(mesh_io_out_c_11_0),
    .io_out_c_11_1(mesh_io_out_c_11_1),
    .io_out_c_12_0(mesh_io_out_c_12_0),
    .io_out_c_12_1(mesh_io_out_c_12_1),
    .io_out_c_13_0(mesh_io_out_c_13_0),
    .io_out_c_13_1(mesh_io_out_c_13_1),
    .io_out_c_14_0(mesh_io_out_c_14_0),
    .io_out_c_14_1(mesh_io_out_c_14_1),
    .io_out_c_15_0(mesh_io_out_c_15_0),
    .io_out_c_15_1(mesh_io_out_c_15_1),
    .io_in_valid_0_0(mesh_io_in_valid_0_0),
    .io_in_valid_0_1(mesh_io_in_valid_0_1),
    .io_in_valid_1_0(mesh_io_in_valid_1_0),
    .io_in_valid_1_1(mesh_io_in_valid_1_1),
    .io_in_valid_2_0(mesh_io_in_valid_2_0),
    .io_in_valid_2_1(mesh_io_in_valid_2_1),
    .io_in_valid_3_0(mesh_io_in_valid_3_0),
    .io_in_valid_3_1(mesh_io_in_valid_3_1),
    .io_in_valid_4_0(mesh_io_in_valid_4_0),
    .io_in_valid_4_1(mesh_io_in_valid_4_1),
    .io_in_valid_5_0(mesh_io_in_valid_5_0),
    .io_in_valid_5_1(mesh_io_in_valid_5_1),
    .io_in_valid_6_0(mesh_io_in_valid_6_0),
    .io_in_valid_6_1(mesh_io_in_valid_6_1),
    .io_in_valid_7_0(mesh_io_in_valid_7_0),
    .io_in_valid_7_1(mesh_io_in_valid_7_1),
    .io_in_valid_8_0(mesh_io_in_valid_8_0),
    .io_in_valid_8_1(mesh_io_in_valid_8_1),
    .io_in_valid_9_0(mesh_io_in_valid_9_0),
    .io_in_valid_9_1(mesh_io_in_valid_9_1),
    .io_in_valid_10_0(mesh_io_in_valid_10_0),
    .io_in_valid_10_1(mesh_io_in_valid_10_1),
    .io_in_valid_11_0(mesh_io_in_valid_11_0),
    .io_in_valid_11_1(mesh_io_in_valid_11_1),
    .io_in_valid_12_0(mesh_io_in_valid_12_0),
    .io_in_valid_12_1(mesh_io_in_valid_12_1),
    .io_in_valid_13_0(mesh_io_in_valid_13_0),
    .io_in_valid_13_1(mesh_io_in_valid_13_1),
    .io_in_valid_14_0(mesh_io_in_valid_14_0),
    .io_in_valid_14_1(mesh_io_in_valid_14_1),
    .io_in_valid_15_0(mesh_io_in_valid_15_0),
    .io_in_valid_15_1(mesh_io_in_valid_15_1),
    .io_out_valid_0_0(mesh_io_out_valid_0_0),
    .io_out_valid_0_1(mesh_io_out_valid_0_1),
    .io_out_valid_1_0(mesh_io_out_valid_1_0),
    .io_out_valid_1_1(mesh_io_out_valid_1_1),
    .io_out_valid_2_0(mesh_io_out_valid_2_0),
    .io_out_valid_2_1(mesh_io_out_valid_2_1),
    .io_out_valid_3_0(mesh_io_out_valid_3_0),
    .io_out_valid_3_1(mesh_io_out_valid_3_1),
    .io_out_valid_4_0(mesh_io_out_valid_4_0),
    .io_out_valid_4_1(mesh_io_out_valid_4_1),
    .io_out_valid_5_0(mesh_io_out_valid_5_0),
    .io_out_valid_5_1(mesh_io_out_valid_5_1),
    .io_out_valid_6_0(mesh_io_out_valid_6_0),
    .io_out_valid_6_1(mesh_io_out_valid_6_1),
    .io_out_valid_7_0(mesh_io_out_valid_7_0),
    .io_out_valid_7_1(mesh_io_out_valid_7_1),
    .io_out_valid_8_0(mesh_io_out_valid_8_0),
    .io_out_valid_8_1(mesh_io_out_valid_8_1),
    .io_out_valid_9_0(mesh_io_out_valid_9_0),
    .io_out_valid_9_1(mesh_io_out_valid_9_1),
    .io_out_valid_10_0(mesh_io_out_valid_10_0),
    .io_out_valid_10_1(mesh_io_out_valid_10_1),
    .io_out_valid_11_0(mesh_io_out_valid_11_0),
    .io_out_valid_11_1(mesh_io_out_valid_11_1),
    .io_out_valid_12_0(mesh_io_out_valid_12_0),
    .io_out_valid_12_1(mesh_io_out_valid_12_1),
    .io_out_valid_13_0(mesh_io_out_valid_13_0),
    .io_out_valid_13_1(mesh_io_out_valid_13_1),
    .io_out_valid_14_0(mesh_io_out_valid_14_0),
    .io_out_valid_14_1(mesh_io_out_valid_14_1),
    .io_out_valid_15_0(mesh_io_out_valid_15_0),
    .io_out_valid_15_1(mesh_io_out_valid_15_1),
    .io_out_control_0_0_dataflow(mesh_io_out_control_0_0_dataflow),
    .io_out_control_0_0_propagate(mesh_io_out_control_0_0_propagate),
    .io_out_control_0_0_shift(mesh_io_out_control_0_0_shift),
    .io_out_control_0_1_dataflow(mesh_io_out_control_0_1_dataflow),
    .io_out_control_0_1_propagate(mesh_io_out_control_0_1_propagate),
    .io_out_control_0_1_shift(mesh_io_out_control_0_1_shift),
    .io_out_control_1_0_dataflow(mesh_io_out_control_1_0_dataflow),
    .io_out_control_1_0_propagate(mesh_io_out_control_1_0_propagate),
    .io_out_control_1_0_shift(mesh_io_out_control_1_0_shift),
    .io_out_control_1_1_dataflow(mesh_io_out_control_1_1_dataflow),
    .io_out_control_1_1_propagate(mesh_io_out_control_1_1_propagate),
    .io_out_control_1_1_shift(mesh_io_out_control_1_1_shift),
    .io_out_control_2_0_dataflow(mesh_io_out_control_2_0_dataflow),
    .io_out_control_2_0_propagate(mesh_io_out_control_2_0_propagate),
    .io_out_control_2_0_shift(mesh_io_out_control_2_0_shift),
    .io_out_control_2_1_dataflow(mesh_io_out_control_2_1_dataflow),
    .io_out_control_2_1_propagate(mesh_io_out_control_2_1_propagate),
    .io_out_control_2_1_shift(mesh_io_out_control_2_1_shift),
    .io_out_control_3_0_dataflow(mesh_io_out_control_3_0_dataflow),
    .io_out_control_3_0_propagate(mesh_io_out_control_3_0_propagate),
    .io_out_control_3_0_shift(mesh_io_out_control_3_0_shift),
    .io_out_control_3_1_dataflow(mesh_io_out_control_3_1_dataflow),
    .io_out_control_3_1_propagate(mesh_io_out_control_3_1_propagate),
    .io_out_control_3_1_shift(mesh_io_out_control_3_1_shift),
    .io_out_control_4_0_dataflow(mesh_io_out_control_4_0_dataflow),
    .io_out_control_4_0_propagate(mesh_io_out_control_4_0_propagate),
    .io_out_control_4_0_shift(mesh_io_out_control_4_0_shift),
    .io_out_control_4_1_dataflow(mesh_io_out_control_4_1_dataflow),
    .io_out_control_4_1_propagate(mesh_io_out_control_4_1_propagate),
    .io_out_control_4_1_shift(mesh_io_out_control_4_1_shift),
    .io_out_control_5_0_dataflow(mesh_io_out_control_5_0_dataflow),
    .io_out_control_5_0_propagate(mesh_io_out_control_5_0_propagate),
    .io_out_control_5_0_shift(mesh_io_out_control_5_0_shift),
    .io_out_control_5_1_dataflow(mesh_io_out_control_5_1_dataflow),
    .io_out_control_5_1_propagate(mesh_io_out_control_5_1_propagate),
    .io_out_control_5_1_shift(mesh_io_out_control_5_1_shift),
    .io_out_control_6_0_dataflow(mesh_io_out_control_6_0_dataflow),
    .io_out_control_6_0_propagate(mesh_io_out_control_6_0_propagate),
    .io_out_control_6_0_shift(mesh_io_out_control_6_0_shift),
    .io_out_control_6_1_dataflow(mesh_io_out_control_6_1_dataflow),
    .io_out_control_6_1_propagate(mesh_io_out_control_6_1_propagate),
    .io_out_control_6_1_shift(mesh_io_out_control_6_1_shift),
    .io_out_control_7_0_dataflow(mesh_io_out_control_7_0_dataflow),
    .io_out_control_7_0_propagate(mesh_io_out_control_7_0_propagate),
    .io_out_control_7_0_shift(mesh_io_out_control_7_0_shift),
    .io_out_control_7_1_dataflow(mesh_io_out_control_7_1_dataflow),
    .io_out_control_7_1_propagate(mesh_io_out_control_7_1_propagate),
    .io_out_control_7_1_shift(mesh_io_out_control_7_1_shift),
    .io_out_control_8_0_dataflow(mesh_io_out_control_8_0_dataflow),
    .io_out_control_8_0_propagate(mesh_io_out_control_8_0_propagate),
    .io_out_control_8_0_shift(mesh_io_out_control_8_0_shift),
    .io_out_control_8_1_dataflow(mesh_io_out_control_8_1_dataflow),
    .io_out_control_8_1_propagate(mesh_io_out_control_8_1_propagate),
    .io_out_control_8_1_shift(mesh_io_out_control_8_1_shift),
    .io_out_control_9_0_dataflow(mesh_io_out_control_9_0_dataflow),
    .io_out_control_9_0_propagate(mesh_io_out_control_9_0_propagate),
    .io_out_control_9_0_shift(mesh_io_out_control_9_0_shift),
    .io_out_control_9_1_dataflow(mesh_io_out_control_9_1_dataflow),
    .io_out_control_9_1_propagate(mesh_io_out_control_9_1_propagate),
    .io_out_control_9_1_shift(mesh_io_out_control_9_1_shift),
    .io_out_control_10_0_dataflow(mesh_io_out_control_10_0_dataflow),
    .io_out_control_10_0_propagate(mesh_io_out_control_10_0_propagate),
    .io_out_control_10_0_shift(mesh_io_out_control_10_0_shift),
    .io_out_control_10_1_dataflow(mesh_io_out_control_10_1_dataflow),
    .io_out_control_10_1_propagate(mesh_io_out_control_10_1_propagate),
    .io_out_control_10_1_shift(mesh_io_out_control_10_1_shift),
    .io_out_control_11_0_dataflow(mesh_io_out_control_11_0_dataflow),
    .io_out_control_11_0_propagate(mesh_io_out_control_11_0_propagate),
    .io_out_control_11_0_shift(mesh_io_out_control_11_0_shift),
    .io_out_control_11_1_dataflow(mesh_io_out_control_11_1_dataflow),
    .io_out_control_11_1_propagate(mesh_io_out_control_11_1_propagate),
    .io_out_control_11_1_shift(mesh_io_out_control_11_1_shift),
    .io_out_control_12_0_dataflow(mesh_io_out_control_12_0_dataflow),
    .io_out_control_12_0_propagate(mesh_io_out_control_12_0_propagate),
    .io_out_control_12_0_shift(mesh_io_out_control_12_0_shift),
    .io_out_control_12_1_dataflow(mesh_io_out_control_12_1_dataflow),
    .io_out_control_12_1_propagate(mesh_io_out_control_12_1_propagate),
    .io_out_control_12_1_shift(mesh_io_out_control_12_1_shift),
    .io_out_control_13_0_dataflow(mesh_io_out_control_13_0_dataflow),
    .io_out_control_13_0_propagate(mesh_io_out_control_13_0_propagate),
    .io_out_control_13_0_shift(mesh_io_out_control_13_0_shift),
    .io_out_control_13_1_dataflow(mesh_io_out_control_13_1_dataflow),
    .io_out_control_13_1_propagate(mesh_io_out_control_13_1_propagate),
    .io_out_control_13_1_shift(mesh_io_out_control_13_1_shift),
    .io_out_control_14_0_dataflow(mesh_io_out_control_14_0_dataflow),
    .io_out_control_14_0_propagate(mesh_io_out_control_14_0_propagate),
    .io_out_control_14_0_shift(mesh_io_out_control_14_0_shift),
    .io_out_control_14_1_dataflow(mesh_io_out_control_14_1_dataflow),
    .io_out_control_14_1_propagate(mesh_io_out_control_14_1_propagate),
    .io_out_control_14_1_shift(mesh_io_out_control_14_1_shift),
    .io_out_control_15_0_dataflow(mesh_io_out_control_15_0_dataflow),
    .io_out_control_15_0_propagate(mesh_io_out_control_15_0_propagate),
    .io_out_control_15_0_shift(mesh_io_out_control_15_0_shift),
    .io_out_control_15_1_dataflow(mesh_io_out_control_15_1_dataflow),
    .io_out_control_15_1_propagate(mesh_io_out_control_15_1_propagate),
    .io_out_control_15_1_shift(mesh_io_out_control_15_1_shift),
    .io_out_id_0_0(mesh_io_out_id_0_0),
    .io_out_id_0_1(mesh_io_out_id_0_1),
    .io_out_id_1_0(mesh_io_out_id_1_0),
    .io_out_id_1_1(mesh_io_out_id_1_1),
    .io_out_id_2_0(mesh_io_out_id_2_0),
    .io_out_id_2_1(mesh_io_out_id_2_1),
    .io_out_id_3_0(mesh_io_out_id_3_0),
    .io_out_id_3_1(mesh_io_out_id_3_1),
    .io_out_id_4_0(mesh_io_out_id_4_0),
    .io_out_id_4_1(mesh_io_out_id_4_1),
    .io_out_id_5_0(mesh_io_out_id_5_0),
    .io_out_id_5_1(mesh_io_out_id_5_1),
    .io_out_id_6_0(mesh_io_out_id_6_0),
    .io_out_id_6_1(mesh_io_out_id_6_1),
    .io_out_id_7_0(mesh_io_out_id_7_0),
    .io_out_id_7_1(mesh_io_out_id_7_1),
    .io_out_id_8_0(mesh_io_out_id_8_0),
    .io_out_id_8_1(mesh_io_out_id_8_1),
    .io_out_id_9_0(mesh_io_out_id_9_0),
    .io_out_id_9_1(mesh_io_out_id_9_1),
    .io_out_id_10_0(mesh_io_out_id_10_0),
    .io_out_id_10_1(mesh_io_out_id_10_1),
    .io_out_id_11_0(mesh_io_out_id_11_0),
    .io_out_id_11_1(mesh_io_out_id_11_1),
    .io_out_id_12_0(mesh_io_out_id_12_0),
    .io_out_id_12_1(mesh_io_out_id_12_1),
    .io_out_id_13_0(mesh_io_out_id_13_0),
    .io_out_id_13_1(mesh_io_out_id_13_1),
    .io_out_id_14_0(mesh_io_out_id_14_0),
    .io_out_id_14_1(mesh_io_out_id_14_1),
    .io_out_id_15_0(mesh_io_out_id_15_0),
    .io_out_id_15_1(mesh_io_out_id_15_1),
    .io_out_last_0_0(mesh_io_out_last_0_0),
    .io_out_last_0_1(mesh_io_out_last_0_1),
    .io_out_last_1_0(mesh_io_out_last_1_0),
    .io_out_last_1_1(mesh_io_out_last_1_1),
    .io_out_last_2_0(mesh_io_out_last_2_0),
    .io_out_last_2_1(mesh_io_out_last_2_1),
    .io_out_last_3_0(mesh_io_out_last_3_0),
    .io_out_last_3_1(mesh_io_out_last_3_1),
    .io_out_last_4_0(mesh_io_out_last_4_0),
    .io_out_last_4_1(mesh_io_out_last_4_1),
    .io_out_last_5_0(mesh_io_out_last_5_0),
    .io_out_last_5_1(mesh_io_out_last_5_1),
    .io_out_last_6_0(mesh_io_out_last_6_0),
    .io_out_last_6_1(mesh_io_out_last_6_1),
    .io_out_last_7_0(mesh_io_out_last_7_0),
    .io_out_last_7_1(mesh_io_out_last_7_1),
    .io_out_last_8_0(mesh_io_out_last_8_0),
    .io_out_last_8_1(mesh_io_out_last_8_1),
    .io_out_last_9_0(mesh_io_out_last_9_0),
    .io_out_last_9_1(mesh_io_out_last_9_1),
    .io_out_last_10_0(mesh_io_out_last_10_0),
    .io_out_last_10_1(mesh_io_out_last_10_1),
    .io_out_last_11_0(mesh_io_out_last_11_0),
    .io_out_last_11_1(mesh_io_out_last_11_1),
    .io_out_last_12_0(mesh_io_out_last_12_0),
    .io_out_last_12_1(mesh_io_out_last_12_1),
    .io_out_last_13_0(mesh_io_out_last_13_0),
    .io_out_last_13_1(mesh_io_out_last_13_1),
    .io_out_last_14_0(mesh_io_out_last_14_0),
    .io_out_last_14_1(mesh_io_out_last_14_1),
    .io_out_last_15_0(mesh_io_out_last_15_0),
    .io_out_last_15_1(mesh_io_out_last_15_1)
  );
  assign io_out_b_0_0 = mesh_io_out_b_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_0_1 = mesh_io_out_b_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_1_0 = mesh_io_out_b_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_1_1 = mesh_io_out_b_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_2_0 = mesh_io_out_b_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_2_1 = mesh_io_out_b_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_3_0 = mesh_io_out_b_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_3_1 = mesh_io_out_b_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_4_0 = mesh_io_out_b_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_4_1 = mesh_io_out_b_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_5_0 = mesh_io_out_b_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_5_1 = mesh_io_out_b_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_6_0 = mesh_io_out_b_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_6_1 = mesh_io_out_b_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_7_0 = mesh_io_out_b_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_7_1 = mesh_io_out_b_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_8_0 = mesh_io_out_b_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_8_1 = mesh_io_out_b_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_9_0 = mesh_io_out_b_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_9_1 = mesh_io_out_b_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_10_0 = mesh_io_out_b_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_10_1 = mesh_io_out_b_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_11_0 = mesh_io_out_b_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_11_1 = mesh_io_out_b_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_12_0 = mesh_io_out_b_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_12_1 = mesh_io_out_b_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_13_0 = mesh_io_out_b_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_13_1 = mesh_io_out_b_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_14_0 = mesh_io_out_b_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_14_1 = mesh_io_out_b_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_15_0 = mesh_io_out_b_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_b_15_1 = mesh_io_out_b_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 69:18]
  assign io_out_c_0_0 = mesh_io_out_c_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_0_1 = mesh_io_out_c_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_1_0 = mesh_io_out_c_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_1_1 = mesh_io_out_c_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_2_0 = mesh_io_out_c_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_2_1 = mesh_io_out_c_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_3_0 = mesh_io_out_c_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_3_1 = mesh_io_out_c_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_4_0 = mesh_io_out_c_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_4_1 = mesh_io_out_c_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_5_0 = mesh_io_out_c_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_5_1 = mesh_io_out_c_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_6_0 = mesh_io_out_c_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_6_1 = mesh_io_out_c_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_7_0 = mesh_io_out_c_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_7_1 = mesh_io_out_c_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_8_0 = mesh_io_out_c_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_8_1 = mesh_io_out_c_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_9_0 = mesh_io_out_c_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_9_1 = mesh_io_out_c_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_10_0 = mesh_io_out_c_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_10_1 = mesh_io_out_c_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_11_0 = mesh_io_out_c_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_11_1 = mesh_io_out_c_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_12_0 = mesh_io_out_c_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_12_1 = mesh_io_out_c_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_13_0 = mesh_io_out_c_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_13_1 = mesh_io_out_c_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_14_0 = mesh_io_out_c_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_14_1 = mesh_io_out_c_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_15_0 = mesh_io_out_c_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_c_15_1 = mesh_io_out_c_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 70:18]
  assign io_out_valid_0_0 = mesh_io_out_valid_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_0_1 = mesh_io_out_valid_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_1_0 = mesh_io_out_valid_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_1_1 = mesh_io_out_valid_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_2_0 = mesh_io_out_valid_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_2_1 = mesh_io_out_valid_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_3_0 = mesh_io_out_valid_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_3_1 = mesh_io_out_valid_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_4_0 = mesh_io_out_valid_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_4_1 = mesh_io_out_valid_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_5_0 = mesh_io_out_valid_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_5_1 = mesh_io_out_valid_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_6_0 = mesh_io_out_valid_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_6_1 = mesh_io_out_valid_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_7_0 = mesh_io_out_valid_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_7_1 = mesh_io_out_valid_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_8_0 = mesh_io_out_valid_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_8_1 = mesh_io_out_valid_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_9_0 = mesh_io_out_valid_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_9_1 = mesh_io_out_valid_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_10_0 = mesh_io_out_valid_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_10_1 = mesh_io_out_valid_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_11_0 = mesh_io_out_valid_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_11_1 = mesh_io_out_valid_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_12_0 = mesh_io_out_valid_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_12_1 = mesh_io_out_valid_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_13_0 = mesh_io_out_valid_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_13_1 = mesh_io_out_valid_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_14_0 = mesh_io_out_valid_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_14_1 = mesh_io_out_valid_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_15_0 = mesh_io_out_valid_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_valid_15_1 = mesh_io_out_valid_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 71:18]
  assign io_out_control_0_0_dataflow = mesh_io_out_control_0_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_0_0_propagate = mesh_io_out_control_0_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_0_0_shift = mesh_io_out_control_0_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_0_1_dataflow = mesh_io_out_control_0_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_0_1_propagate = mesh_io_out_control_0_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_0_1_shift = mesh_io_out_control_0_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_1_0_dataflow = mesh_io_out_control_1_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_1_0_propagate = mesh_io_out_control_1_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_1_0_shift = mesh_io_out_control_1_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_1_1_dataflow = mesh_io_out_control_1_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_1_1_propagate = mesh_io_out_control_1_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_1_1_shift = mesh_io_out_control_1_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_2_0_dataflow = mesh_io_out_control_2_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_2_0_propagate = mesh_io_out_control_2_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_2_0_shift = mesh_io_out_control_2_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_2_1_dataflow = mesh_io_out_control_2_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_2_1_propagate = mesh_io_out_control_2_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_2_1_shift = mesh_io_out_control_2_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_3_0_dataflow = mesh_io_out_control_3_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_3_0_propagate = mesh_io_out_control_3_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_3_0_shift = mesh_io_out_control_3_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_3_1_dataflow = mesh_io_out_control_3_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_3_1_propagate = mesh_io_out_control_3_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_3_1_shift = mesh_io_out_control_3_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_4_0_dataflow = mesh_io_out_control_4_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_4_0_propagate = mesh_io_out_control_4_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_4_0_shift = mesh_io_out_control_4_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_4_1_dataflow = mesh_io_out_control_4_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_4_1_propagate = mesh_io_out_control_4_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_4_1_shift = mesh_io_out_control_4_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_5_0_dataflow = mesh_io_out_control_5_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_5_0_propagate = mesh_io_out_control_5_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_5_0_shift = mesh_io_out_control_5_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_5_1_dataflow = mesh_io_out_control_5_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_5_1_propagate = mesh_io_out_control_5_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_5_1_shift = mesh_io_out_control_5_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_6_0_dataflow = mesh_io_out_control_6_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_6_0_propagate = mesh_io_out_control_6_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_6_0_shift = mesh_io_out_control_6_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_6_1_dataflow = mesh_io_out_control_6_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_6_1_propagate = mesh_io_out_control_6_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_6_1_shift = mesh_io_out_control_6_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_7_0_dataflow = mesh_io_out_control_7_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_7_0_propagate = mesh_io_out_control_7_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_7_0_shift = mesh_io_out_control_7_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_7_1_dataflow = mesh_io_out_control_7_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_7_1_propagate = mesh_io_out_control_7_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_7_1_shift = mesh_io_out_control_7_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_8_0_dataflow = mesh_io_out_control_8_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_8_0_propagate = mesh_io_out_control_8_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_8_0_shift = mesh_io_out_control_8_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_8_1_dataflow = mesh_io_out_control_8_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_8_1_propagate = mesh_io_out_control_8_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_8_1_shift = mesh_io_out_control_8_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_9_0_dataflow = mesh_io_out_control_9_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_9_0_propagate = mesh_io_out_control_9_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_9_0_shift = mesh_io_out_control_9_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_9_1_dataflow = mesh_io_out_control_9_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_9_1_propagate = mesh_io_out_control_9_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_9_1_shift = mesh_io_out_control_9_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_10_0_dataflow = mesh_io_out_control_10_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_10_0_propagate = mesh_io_out_control_10_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_10_0_shift = mesh_io_out_control_10_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_10_1_dataflow = mesh_io_out_control_10_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_10_1_propagate = mesh_io_out_control_10_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_10_1_shift = mesh_io_out_control_10_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_11_0_dataflow = mesh_io_out_control_11_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_11_0_propagate = mesh_io_out_control_11_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_11_0_shift = mesh_io_out_control_11_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_11_1_dataflow = mesh_io_out_control_11_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_11_1_propagate = mesh_io_out_control_11_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_11_1_shift = mesh_io_out_control_11_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_12_0_dataflow = mesh_io_out_control_12_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_12_0_propagate = mesh_io_out_control_12_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_12_0_shift = mesh_io_out_control_12_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_12_1_dataflow = mesh_io_out_control_12_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_12_1_propagate = mesh_io_out_control_12_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_12_1_shift = mesh_io_out_control_12_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_13_0_dataflow = mesh_io_out_control_13_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_13_0_propagate = mesh_io_out_control_13_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_13_0_shift = mesh_io_out_control_13_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_13_1_dataflow = mesh_io_out_control_13_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_13_1_propagate = mesh_io_out_control_13_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_13_1_shift = mesh_io_out_control_13_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_14_0_dataflow = mesh_io_out_control_14_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_14_0_propagate = mesh_io_out_control_14_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_14_0_shift = mesh_io_out_control_14_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_14_1_dataflow = mesh_io_out_control_14_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_14_1_propagate = mesh_io_out_control_14_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_14_1_shift = mesh_io_out_control_14_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_15_0_dataflow = mesh_io_out_control_15_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_15_0_propagate = mesh_io_out_control_15_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_15_0_shift = mesh_io_out_control_15_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_15_1_dataflow = mesh_io_out_control_15_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_15_1_propagate = mesh_io_out_control_15_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_control_15_1_shift = mesh_io_out_control_15_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 72:18]
  assign io_out_id_0_0 = mesh_io_out_id_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_0_1 = mesh_io_out_id_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_1_0 = mesh_io_out_id_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_1_1 = mesh_io_out_id_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_2_0 = mesh_io_out_id_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_2_1 = mesh_io_out_id_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_3_0 = mesh_io_out_id_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_3_1 = mesh_io_out_id_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_4_0 = mesh_io_out_id_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_4_1 = mesh_io_out_id_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_5_0 = mesh_io_out_id_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_5_1 = mesh_io_out_id_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_6_0 = mesh_io_out_id_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_6_1 = mesh_io_out_id_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_7_0 = mesh_io_out_id_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_7_1 = mesh_io_out_id_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_8_0 = mesh_io_out_id_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_8_1 = mesh_io_out_id_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_9_0 = mesh_io_out_id_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_9_1 = mesh_io_out_id_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_10_0 = mesh_io_out_id_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_10_1 = mesh_io_out_id_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_11_0 = mesh_io_out_id_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_11_1 = mesh_io_out_id_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_12_0 = mesh_io_out_id_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_12_1 = mesh_io_out_id_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_13_0 = mesh_io_out_id_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_13_1 = mesh_io_out_id_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_14_0 = mesh_io_out_id_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_14_1 = mesh_io_out_id_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_15_0 = mesh_io_out_id_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_id_15_1 = mesh_io_out_id_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 73:18]
  assign io_out_last_0_0 = mesh_io_out_last_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_0_1 = mesh_io_out_last_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_1_0 = mesh_io_out_last_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_1_1 = mesh_io_out_last_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_2_0 = mesh_io_out_last_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_2_1 = mesh_io_out_last_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_3_0 = mesh_io_out_last_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_3_1 = mesh_io_out_last_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_4_0 = mesh_io_out_last_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_4_1 = mesh_io_out_last_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_5_0 = mesh_io_out_last_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_5_1 = mesh_io_out_last_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_6_0 = mesh_io_out_last_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_6_1 = mesh_io_out_last_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_7_0 = mesh_io_out_last_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_7_1 = mesh_io_out_last_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_8_0 = mesh_io_out_last_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_8_1 = mesh_io_out_last_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_9_0 = mesh_io_out_last_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_9_1 = mesh_io_out_last_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_10_0 = mesh_io_out_last_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_10_1 = mesh_io_out_last_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_11_0 = mesh_io_out_last_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_11_1 = mesh_io_out_last_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_12_0 = mesh_io_out_last_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_12_1 = mesh_io_out_last_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_13_0 = mesh_io_out_last_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_13_1 = mesh_io_out_last_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_14_0 = mesh_io_out_last_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_14_1 = mesh_io_out_last_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_15_0 = mesh_io_out_last_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign io_out_last_15_1 = mesh_io_out_last_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 74:18]
  assign mesh_clock = clock;
  assign mesh_io_in_a_0_0 = io_in_a_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_0_1 = io_in_a_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_1_0 = io_in_a_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_1_1 = io_in_a_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_2_0 = io_in_a_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_2_1 = io_in_a_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_3_0 = io_in_a_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_3_1 = io_in_a_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_4_0 = io_in_a_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_4_1 = io_in_a_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_5_0 = io_in_a_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_5_1 = io_in_a_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_6_0 = io_in_a_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_6_1 = io_in_a_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_7_0 = io_in_a_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_7_1 = io_in_a_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_8_0 = io_in_a_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_8_1 = io_in_a_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_9_0 = io_in_a_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_9_1 = io_in_a_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_10_0 = io_in_a_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_10_1 = io_in_a_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_11_0 = io_in_a_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_11_1 = io_in_a_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_12_0 = io_in_a_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_12_1 = io_in_a_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_13_0 = io_in_a_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_13_1 = io_in_a_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_14_0 = io_in_a_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_14_1 = io_in_a_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_15_0 = io_in_a_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_a_15_1 = io_in_a_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 60:22]
  assign mesh_io_in_b_0_0 = io_in_b_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_0_1 = io_in_b_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_1_0 = io_in_b_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_1_1 = io_in_b_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_2_0 = io_in_b_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_2_1 = io_in_b_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_3_0 = io_in_b_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_3_1 = io_in_b_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_4_0 = io_in_b_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_4_1 = io_in_b_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_5_0 = io_in_b_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_5_1 = io_in_b_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_6_0 = io_in_b_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_6_1 = io_in_b_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_7_0 = io_in_b_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_7_1 = io_in_b_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_8_0 = io_in_b_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_8_1 = io_in_b_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_9_0 = io_in_b_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_9_1 = io_in_b_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_10_0 = io_in_b_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_10_1 = io_in_b_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_11_0 = io_in_b_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_11_1 = io_in_b_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_12_0 = io_in_b_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_12_1 = io_in_b_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_13_0 = io_in_b_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_13_1 = io_in_b_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_14_0 = io_in_b_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_14_1 = io_in_b_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_15_0 = io_in_b_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_b_15_1 = io_in_b_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 61:22]
  assign mesh_io_in_d_0_0 = io_in_d_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_0_1 = io_in_d_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_1_0 = io_in_d_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_1_1 = io_in_d_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_2_0 = io_in_d_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_2_1 = io_in_d_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_3_0 = io_in_d_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_3_1 = io_in_d_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_4_0 = io_in_d_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_4_1 = io_in_d_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_5_0 = io_in_d_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_5_1 = io_in_d_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_6_0 = io_in_d_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_6_1 = io_in_d_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_7_0 = io_in_d_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_7_1 = io_in_d_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_8_0 = io_in_d_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_8_1 = io_in_d_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_9_0 = io_in_d_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_9_1 = io_in_d_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_10_0 = io_in_d_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_10_1 = io_in_d_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_11_0 = io_in_d_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_11_1 = io_in_d_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_12_0 = io_in_d_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_12_1 = io_in_d_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_13_0 = io_in_d_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_13_1 = io_in_d_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_14_0 = io_in_d_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_14_1 = io_in_d_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_15_0 = io_in_d_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_d_15_1 = io_in_d_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 62:22]
  assign mesh_io_in_control_0_0_dataflow = io_in_control_0_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_0_0_propagate = io_in_control_0_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_0_0_shift = io_in_control_0_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_0_1_dataflow = io_in_control_0_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_0_1_propagate = io_in_control_0_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_0_1_shift = io_in_control_0_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_1_0_dataflow = io_in_control_1_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_1_0_propagate = io_in_control_1_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_1_0_shift = io_in_control_1_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_1_1_dataflow = io_in_control_1_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_1_1_propagate = io_in_control_1_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_1_1_shift = io_in_control_1_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_2_0_dataflow = io_in_control_2_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_2_0_propagate = io_in_control_2_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_2_0_shift = io_in_control_2_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_2_1_dataflow = io_in_control_2_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_2_1_propagate = io_in_control_2_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_2_1_shift = io_in_control_2_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_3_0_dataflow = io_in_control_3_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_3_0_propagate = io_in_control_3_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_3_0_shift = io_in_control_3_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_3_1_dataflow = io_in_control_3_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_3_1_propagate = io_in_control_3_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_3_1_shift = io_in_control_3_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_4_0_dataflow = io_in_control_4_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_4_0_propagate = io_in_control_4_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_4_0_shift = io_in_control_4_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_4_1_dataflow = io_in_control_4_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_4_1_propagate = io_in_control_4_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_4_1_shift = io_in_control_4_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_5_0_dataflow = io_in_control_5_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_5_0_propagate = io_in_control_5_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_5_0_shift = io_in_control_5_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_5_1_dataflow = io_in_control_5_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_5_1_propagate = io_in_control_5_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_5_1_shift = io_in_control_5_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_6_0_dataflow = io_in_control_6_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_6_0_propagate = io_in_control_6_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_6_0_shift = io_in_control_6_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_6_1_dataflow = io_in_control_6_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_6_1_propagate = io_in_control_6_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_6_1_shift = io_in_control_6_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_7_0_dataflow = io_in_control_7_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_7_0_propagate = io_in_control_7_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_7_0_shift = io_in_control_7_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_7_1_dataflow = io_in_control_7_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_7_1_propagate = io_in_control_7_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_7_1_shift = io_in_control_7_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_8_0_dataflow = io_in_control_8_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_8_0_propagate = io_in_control_8_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_8_0_shift = io_in_control_8_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_8_1_dataflow = io_in_control_8_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_8_1_propagate = io_in_control_8_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_8_1_shift = io_in_control_8_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_9_0_dataflow = io_in_control_9_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_9_0_propagate = io_in_control_9_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_9_0_shift = io_in_control_9_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_9_1_dataflow = io_in_control_9_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_9_1_propagate = io_in_control_9_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_9_1_shift = io_in_control_9_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_10_0_dataflow = io_in_control_10_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_10_0_propagate = io_in_control_10_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_10_0_shift = io_in_control_10_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_10_1_dataflow = io_in_control_10_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_10_1_propagate = io_in_control_10_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_10_1_shift = io_in_control_10_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_11_0_dataflow = io_in_control_11_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_11_0_propagate = io_in_control_11_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_11_0_shift = io_in_control_11_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_11_1_dataflow = io_in_control_11_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_11_1_propagate = io_in_control_11_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_11_1_shift = io_in_control_11_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_12_0_dataflow = io_in_control_12_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_12_0_propagate = io_in_control_12_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_12_0_shift = io_in_control_12_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_12_1_dataflow = io_in_control_12_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_12_1_propagate = io_in_control_12_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_12_1_shift = io_in_control_12_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_13_0_dataflow = io_in_control_13_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_13_0_propagate = io_in_control_13_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_13_0_shift = io_in_control_13_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_13_1_dataflow = io_in_control_13_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_13_1_propagate = io_in_control_13_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_13_1_shift = io_in_control_13_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_14_0_dataflow = io_in_control_14_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_14_0_propagate = io_in_control_14_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_14_0_shift = io_in_control_14_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_14_1_dataflow = io_in_control_14_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_14_1_propagate = io_in_control_14_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_14_1_shift = io_in_control_14_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_15_0_dataflow = io_in_control_15_0_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_15_0_propagate = io_in_control_15_0_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_15_0_shift = io_in_control_15_0_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_15_1_dataflow = io_in_control_15_1_dataflow; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_15_1_propagate = io_in_control_15_1_propagate; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_control_15_1_shift = io_in_control_15_1_shift; // @[src/main/scala/gemmini/GemminiMeshTop.scala 63:22]
  assign mesh_io_in_id_0_0 = io_in_id_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_0_1 = io_in_id_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_1_0 = io_in_id_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_1_1 = io_in_id_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_2_0 = io_in_id_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_2_1 = io_in_id_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_3_0 = io_in_id_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_3_1 = io_in_id_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_4_0 = io_in_id_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_4_1 = io_in_id_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_5_0 = io_in_id_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_5_1 = io_in_id_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_6_0 = io_in_id_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_6_1 = io_in_id_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_7_0 = io_in_id_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_7_1 = io_in_id_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_8_0 = io_in_id_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_8_1 = io_in_id_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_9_0 = io_in_id_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_9_1 = io_in_id_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_10_0 = io_in_id_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_10_1 = io_in_id_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_11_0 = io_in_id_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_11_1 = io_in_id_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_12_0 = io_in_id_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_12_1 = io_in_id_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_13_0 = io_in_id_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_13_1 = io_in_id_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_14_0 = io_in_id_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_14_1 = io_in_id_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_15_0 = io_in_id_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_id_15_1 = io_in_id_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 64:22]
  assign mesh_io_in_last_0_0 = io_in_last_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_0_1 = io_in_last_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_1_0 = io_in_last_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_1_1 = io_in_last_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_2_0 = io_in_last_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_2_1 = io_in_last_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_3_0 = io_in_last_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_3_1 = io_in_last_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_4_0 = io_in_last_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_4_1 = io_in_last_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_5_0 = io_in_last_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_5_1 = io_in_last_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_6_0 = io_in_last_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_6_1 = io_in_last_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_7_0 = io_in_last_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_7_1 = io_in_last_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_8_0 = io_in_last_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_8_1 = io_in_last_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_9_0 = io_in_last_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_9_1 = io_in_last_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_10_0 = io_in_last_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_10_1 = io_in_last_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_11_0 = io_in_last_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_11_1 = io_in_last_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_12_0 = io_in_last_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_12_1 = io_in_last_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_13_0 = io_in_last_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_13_1 = io_in_last_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_14_0 = io_in_last_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_14_1 = io_in_last_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_15_0 = io_in_last_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_last_15_1 = io_in_last_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 65:22]
  assign mesh_io_in_valid_0_0 = io_in_valid_0_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_0_1 = io_in_valid_0_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_1_0 = io_in_valid_1_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_1_1 = io_in_valid_1_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_2_0 = io_in_valid_2_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_2_1 = io_in_valid_2_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_3_0 = io_in_valid_3_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_3_1 = io_in_valid_3_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_4_0 = io_in_valid_4_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_4_1 = io_in_valid_4_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_5_0 = io_in_valid_5_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_5_1 = io_in_valid_5_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_6_0 = io_in_valid_6_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_6_1 = io_in_valid_6_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_7_0 = io_in_valid_7_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_7_1 = io_in_valid_7_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_8_0 = io_in_valid_8_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_8_1 = io_in_valid_8_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_9_0 = io_in_valid_9_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_9_1 = io_in_valid_9_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_10_0 = io_in_valid_10_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_10_1 = io_in_valid_10_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_11_0 = io_in_valid_11_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_11_1 = io_in_valid_11_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_12_0 = io_in_valid_12_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_12_1 = io_in_valid_12_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_13_0 = io_in_valid_13_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_13_1 = io_in_valid_13_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_14_0 = io_in_valid_14_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_14_1 = io_in_valid_14_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_15_0 = io_in_valid_15_0; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
  assign mesh_io_in_valid_15_1 = io_in_valid_15_1; // @[src/main/scala/gemmini/GemminiMeshTop.scala 66:22]
endmodule
